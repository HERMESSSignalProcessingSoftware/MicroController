-- Version: v12.6 12.900.20.24
-- File used only for Simulation

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sdf_IOPAD_TRI is

    port( PAD : out   std_logic;
          D   : in    std_logic;
          E   : in    std_logic
        );

end sdf_IOPAD_TRI;

architecture DEF_ARCH of sdf_IOPAD_TRI is 

  component IOPAD_TRI_VDDI
    port( OIN_VDD : in    std_logic := 'U';
          EIN_VDD : in    std_logic := 'U';
          PAD_P   : out   std_logic
        );
  end component;

  component IOPAD_VDD
    port( OIN_P    : in    std_logic := 'U';
          EIN_P    : in    std_logic := 'U';
          IOUT_VDD : in    std_logic := 'U';
          OIN_VDD  : out   std_logic;
          EIN_VDD  : out   std_logic;
          IOUT_IN  : out   std_logic
        );
  end component;

    signal NET_OIN_VDD, NET_EIN_VDD : std_logic;

begin 


    U_VCCI : IOPAD_TRI_VDDI
      port map(OIN_VDD => NET_OIN_VDD, EIN_VDD => NET_EIN_VDD, 
        PAD_P => PAD);
    
    U_VCCA : IOPAD_VDD
      port map(OIN_P => D, EIN_P => E, IOUT_VDD => OPEN, OIN_VDD
         => NET_OIN_VDD, EIN_VDD => NET_EIN_VDD, IOUT_IN => OPEN);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sdf_IOPAD_IN is

    port( PAD : in    std_logic;
          Y   : out   std_logic
        );

end sdf_IOPAD_IN;

architecture DEF_ARCH of sdf_IOPAD_IN is 

  component IOPAD_IN_VDDI
    port( PAD_P    : in    std_logic := 'U';
          IOUT_VDD : out   std_logic
        );
  end component;

  component IOPAD_DELAY
    port( IOUT_IN : in    std_logic := 'U';
          IOUT_P  : out   std_logic
        );
  end component;

  component IOPAD_VDD
    port( OIN_P    : in    std_logic := 'U';
          EIN_P    : in    std_logic := 'U';
          IOUT_VDD : in    std_logic := 'U';
          OIN_VDD  : out   std_logic;
          EIN_VDD  : out   std_logic;
          IOUT_IN  : out   std_logic
        );
  end component;

  component GND
    port(Y : out std_logic); 
  end component;

    signal NET_IOUT_VDD, NET_IOUT_IN, ADLIB_GND : std_logic;
    signal GND_power_net1 : std_logic;

begin 

    ADLIB_GND <= GND_power_net1;

    U_VCCI : IOPAD_IN_VDDI
      port map(PAD_P => PAD, IOUT_VDD => NET_IOUT_VDD);
    
    U_DELAY : IOPAD_DELAY
      port map(IOUT_IN => NET_IOUT_IN, IOUT_P => Y);
    
    U_VCCA : IOPAD_VDD
      port map(OIN_P => ADLIB_GND, EIN_P => ADLIB_GND, IOUT_VDD
         => NET_IOUT_VDD, OIN_VDD => OPEN, EIN_VDD => OPEN, 
        IOUT_IN => NET_IOUT_IN);
    
    GND_power_inst1 : GND
      port map( Y => GND_power_net1);


end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sb is

    port( DEVRST_N           : in    std_logic;
          MISO               : in    std_logic;
          MMUART_0_RXD_F2M   : in    std_logic;
          RXSM_LO            : in    std_logic;
          RXSM_SODS          : in    std_logic;
          RXSM_SOE           : in    std_logic;
          stamp0_ready_dms1  : in    std_logic;
          stamp0_ready_dms2  : in    std_logic;
          stamp0_ready_temp  : in    std_logic;
          stamp0_spi_miso    : in    std_logic;
          ENABLE_MEMORY_LED  : out   std_logic;
          LED_HEARTBEAT      : out   std_logic;
          LED_RECORDING      : out   std_logic;
          MMUART_0_TXD_M2F   : out   std_logic;
          MOSI               : out   std_logic;
          SCLK               : out   std_logic;
          adc_clk            : out   std_logic;
          adc_start          : out   std_logic;
          debug_led          : out   std_logic;
          nCS1               : out   std_logic;
          nCS2               : out   std_logic;
          resetn             : out   std_logic;
          stamp0_spi_clock   : out   std_logic;
          stamp0_spi_dms1_cs : out   std_logic;
          stamp0_spi_dms2_cs : out   std_logic;
          stamp0_spi_mosi    : out   std_logic;
          stamp0_spi_temp_cs : out   std_logic
        );

end sb;

architecture DEF_ARCH of sb is 

  component IP_INTERFACE
    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          IPA : out   std_logic;
          IPB : out   std_logic;
          IPC : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1_CC
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic;
          CC  : in    std_logic := 'U';
          P   : out   std_logic;
          UB  : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV_BA
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RGB_NG
    port( An  : in    std_logic := 'U';
          ENn : in    std_logic := 'U';
          YL  : out   std_logic;
          YR  : out   std_logic
        );
  end component;

  component sdf_IOPAD_TRI
    port( PAD : out   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U'
        );
  end component;

  component CC_CONFIG
    port( CI : in    std_logic := 'U';
          CO : out   std_logic;
          P  : in    std_logic_vector(0 to 11) := (others => 'U');
          UB : in    std_logic_vector(0 to 11) := (others => 'U');
          CC : out   std_logic_vector(0 to 11)
        );
  end component;

  component GB_NG
    port( An  : in    std_logic := 'U';
          ENn : in    std_logic := 'U';
          YNn : out   std_logic;
          YSn : out   std_logic
        );
  end component;

  component IOTRI_OB_EB
    port( D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          DOUT : out   std_logic;
          EOUT : out   std_logic
        );
  end component;

  component IOENFF_BYPASS
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOINFF_BYPASS
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOIN_IB
    port( YIN : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component sdf_IOPAD_IN
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component IOOUTFF_BYPASS
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

  component FCEND_BUFF_CC
    port( FCI : in    std_logic := 'U';
          CO  : out   std_logic;
          CC  : in    std_logic := 'U';
          P   : out   std_logic;
          UB  : out   std_logic
        );
  end component;

  component CFG0
    generic (INIT:std_logic_vector(0 downto 0) := "0");

    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MSS_010_IP

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic
        );
  end component;

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component SYSRESET_FF
    port( UDRCAP           : out   std_logic;
          UDRSH            : out   std_logic;
          UDRUPD           : out   std_logic;
          UIREG            : out   std_logic_vector(7 downto 0);
          URSTB            : out   std_logic;
          UDRCK            : out   std_logic;
          UTDI             : out   std_logic;
          POWER_ON_RESET_N : out   std_logic;
          FF_TO_START      : out   std_logic;
          FF_DONE          : out   std_logic;
          UTDO             : in    std_logic := 'U';
          DEVRST_N         : in    std_logic := 'U';
          TDI              : in    std_logic := 'U';
          TMS              : in    std_logic := 'U';
          TCK              : in    std_logic := 'U';
          TRSTB            : in    std_logic := 'U';
          TDO              : out   std_logic
        );
  end component;

  component GND
    port(Y : out std_logic); 
  end component;

  component VCC
    port(Y : out std_logic); 
  end component;

    signal \sb_sb_0_STAMP_PADDR[11]\, \sb_sb_0_STAMP_PADDR[10]\, 
        \sb_sb_0_STAMP_PADDR[9]\, \sb_sb_0_STAMP_PADDR[8]\, 
        \sb_sb_0_STAMP_PADDR[7]\, \sb_sb_0_STAMP_PADDR[6]\, 
        \sb_sb_0_STAMP_PADDR[5]\, \sb_sb_0_STAMP_PADDR[4]\, 
        \sb_sb_0_STAMP_PADDR[3]\, \sb_sb_0_STAMP_PADDR[2]\, 
        \sb_sb_0_STAMP_PADDR[1]\, \sb_sb_0_STAMP_PADDR[0]\, 
        \sb_sb_0_Memory_PRDATA[31]\, \sb_sb_0_Memory_PRDATA[30]\, 
        \sb_sb_0_Memory_PRDATA[29]\, \sb_sb_0_Memory_PRDATA[28]\, 
        \sb_sb_0_Memory_PRDATA[27]\, \sb_sb_0_Memory_PRDATA[26]\, 
        \sb_sb_0_Memory_PRDATA[25]\, \sb_sb_0_Memory_PRDATA[24]\, 
        \sb_sb_0_Memory_PRDATA[23]\, \sb_sb_0_Memory_PRDATA[22]\, 
        \sb_sb_0_Memory_PRDATA[21]\, \sb_sb_0_Memory_PRDATA[20]\, 
        \sb_sb_0_Memory_PRDATA[19]\, \sb_sb_0_Memory_PRDATA[18]\, 
        \sb_sb_0_Memory_PRDATA[17]\, \sb_sb_0_Memory_PRDATA[16]\, 
        \sb_sb_0_Memory_PRDATA[15]\, \sb_sb_0_Memory_PRDATA[14]\, 
        \sb_sb_0_Memory_PRDATA[13]\, \sb_sb_0_Memory_PRDATA[12]\, 
        \sb_sb_0_Memory_PRDATA[11]\, \sb_sb_0_Memory_PRDATA[10]\, 
        \sb_sb_0_Memory_PRDATA[9]\, \sb_sb_0_Memory_PRDATA[8]\, 
        \sb_sb_0_Memory_PRDATA[7]\, \sb_sb_0_Memory_PRDATA[6]\, 
        \sb_sb_0_Memory_PRDATA[5]\, \sb_sb_0_Memory_PRDATA[4]\, 
        \sb_sb_0_Memory_PRDATA[3]\, \sb_sb_0_Memory_PRDATA[2]\, 
        \sb_sb_0_Memory_PRDATA[1]\, \sb_sb_0_Memory_PRDATA[0]\, 
        \sb_sb_0_STAMP_PRDATA[31]\, \sb_sb_0_STAMP_PRDATA[30]\, 
        \sb_sb_0_STAMP_PRDATA[29]\, \sb_sb_0_STAMP_PRDATA[28]\, 
        \sb_sb_0_STAMP_PRDATA[27]\, \sb_sb_0_STAMP_PRDATA[26]\, 
        \sb_sb_0_STAMP_PRDATA[25]\, \sb_sb_0_STAMP_PRDATA[24]\, 
        \sb_sb_0_STAMP_PRDATA[23]\, \sb_sb_0_STAMP_PRDATA[22]\, 
        \sb_sb_0_STAMP_PRDATA[21]\, \sb_sb_0_STAMP_PRDATA[20]\, 
        \sb_sb_0_STAMP_PRDATA[19]\, \sb_sb_0_STAMP_PRDATA[18]\, 
        \sb_sb_0_STAMP_PRDATA[17]\, \sb_sb_0_STAMP_PRDATA[16]\, 
        \sb_sb_0_STAMP_PRDATA[15]\, \sb_sb_0_STAMP_PRDATA[14]\, 
        \sb_sb_0_STAMP_PRDATA[13]\, \sb_sb_0_STAMP_PRDATA[12]\, 
        \sb_sb_0_STAMP_PRDATA[11]\, \sb_sb_0_STAMP_PRDATA[10]\, 
        \sb_sb_0_STAMP_PRDATA[9]\, \sb_sb_0_STAMP_PRDATA[8]\, 
        \sb_sb_0_STAMP_PRDATA[7]\, \sb_sb_0_STAMP_PRDATA[6]\, 
        \sb_sb_0_STAMP_PRDATA[5]\, \sb_sb_0_STAMP_PRDATA[4]\, 
        \sb_sb_0_STAMP_PRDATA[3]\, \sb_sb_0_STAMP_PRDATA[2]\, 
        \sb_sb_0_STAMP_PRDATA[1]\, \sb_sb_0_STAMP_PRDATA[0]\, 
        \STAMP_0_data_frame[63]\, \STAMP_0_data_frame[62]\, 
        \STAMP_0_data_frame[61]\, \STAMP_0_data_frame[60]\, 
        \STAMP_0_data_frame[59]\, \STAMP_0_data_frame[58]\, 
        \STAMP_0_data_frame[57]\, \STAMP_0_data_frame[56]\, 
        \STAMP_0_data_frame[55]\, \STAMP_0_data_frame[54]\, 
        \STAMP_0_data_frame[53]\, \STAMP_0_data_frame[52]\, 
        \STAMP_0_data_frame[51]\, \STAMP_0_data_frame[50]\, 
        \STAMP_0_data_frame[49]\, \STAMP_0_data_frame[48]\, 
        \STAMP_0_data_frame[47]\, \STAMP_0_data_frame[46]\, 
        \STAMP_0_data_frame[45]\, \STAMP_0_data_frame[44]\, 
        \STAMP_0_data_frame[43]\, \STAMP_0_data_frame[42]\, 
        \STAMP_0_data_frame[41]\, \STAMP_0_data_frame[40]\, 
        \STAMP_0_data_frame[39]\, \STAMP_0_data_frame[38]\, 
        \STAMP_0_data_frame[37]\, \STAMP_0_data_frame[36]\, 
        \STAMP_0_data_frame[35]\, \STAMP_0_data_frame[34]\, 
        \STAMP_0_data_frame[33]\, \STAMP_0_data_frame[32]\, 
        \STAMP_0_data_frame[31]\, \STAMP_0_data_frame[30]\, 
        \STAMP_0_data_frame[29]\, \STAMP_0_data_frame[28]\, 
        \STAMP_0_data_frame[27]\, \STAMP_0_data_frame[26]\, 
        \STAMP_0_data_frame[25]\, \STAMP_0_data_frame[24]\, 
        \STAMP_0_data_frame[23]\, \STAMP_0_data_frame[22]\, 
        \STAMP_0_data_frame[21]\, \STAMP_0_data_frame[20]\, 
        \STAMP_0_data_frame[19]\, \STAMP_0_data_frame[18]\, 
        \STAMP_0_data_frame[17]\, \STAMP_0_data_frame[16]\, 
        \STAMP_0_data_frame[15]\, \STAMP_0_data_frame[14]\, 
        \STAMP_0_data_frame[13]\, \STAMP_0_data_frame[12]\, 
        \STAMP_0_data_frame[11]\, \STAMP_0_data_frame[10]\, 
        \STAMP_0_data_frame[9]\, \STAMP_0_data_frame[8]\, 
        \STAMP_0_data_frame[7]\, \STAMP_0_data_frame[6]\, 
        \STAMP_0_data_frame[5]\, \STAMP_0_data_frame[4]\, 
        \STAMP_0_data_frame[3]\, \STAMP_0_data_frame[2]\, 
        \STAMP_0_data_frame[1]\, \STAMP_0_data_frame[0]\, 
        \sb_sb_0_STAMP_PWDATA[31]\, \sb_sb_0_STAMP_PWDATA[30]\, 
        \sb_sb_0_STAMP_PWDATA[29]\, \sb_sb_0_STAMP_PWDATA[28]\, 
        \sb_sb_0_STAMP_PWDATA[27]\, \sb_sb_0_STAMP_PWDATA[26]\, 
        \sb_sb_0_STAMP_PWDATA[25]\, \sb_sb_0_STAMP_PWDATA[24]\, 
        \sb_sb_0_STAMP_PWDATA[23]\, \sb_sb_0_STAMP_PWDATA[22]\, 
        \sb_sb_0_STAMP_PWDATA[21]\, \sb_sb_0_STAMP_PWDATA[20]\, 
        \sb_sb_0_STAMP_PWDATA[19]\, \sb_sb_0_STAMP_PWDATA[18]\, 
        \sb_sb_0_STAMP_PWDATA[17]\, \sb_sb_0_STAMP_PWDATA[16]\, 
        \sb_sb_0_STAMP_PWDATA[15]\, \sb_sb_0_STAMP_PWDATA[14]\, 
        \sb_sb_0_STAMP_PWDATA[13]\, \sb_sb_0_STAMP_PWDATA[12]\, 
        \sb_sb_0_STAMP_PWDATA[11]\, \sb_sb_0_STAMP_PWDATA[10]\, 
        \sb_sb_0_STAMP_PWDATA[9]\, \sb_sb_0_STAMP_PWDATA[8]\, 
        \sb_sb_0_STAMP_PWDATA[7]\, \sb_sb_0_STAMP_PWDATA[6]\, 
        \sb_sb_0_STAMP_PWDATA[5]\, \sb_sb_0_STAMP_PWDATA[4]\, 
        \sb_sb_0_STAMP_PWDATA[3]\, \sb_sb_0_STAMP_PWDATA[2]\, 
        \sb_sb_0_STAMP_PWDATA[1]\, \sb_sb_0_STAMP_PWDATA[0]\, 
        sb_sb_0_GPIO_3_M2F, \sb_sb_0/CCC_0/GL0_INST/U0_YNn\, 
        STAMP_0_new_avail, MemorySynchronizer_0_dataReadyReset, 
        MemorySynchronizer_0_SynchronizerInterrupt, 
        MemorySynchronizer_0_ReadInterrupt, sb_sb_0_Memory_PSELx, 
        sb_sb_0_STAMP_PENABLE, sb_sb_0_STAMP_PWRITE, 
        sb_sb_0_Memory_PREADY, sb_sb_0_POWER_ON_RESET_N, 
        sb_sb_0_GPIO_4_M2F, sb_sb_0_STAMP_PREADY, mosi_1, 
        \AND2_0_RNIKOS1/U0_YNn\, NN_1, debug_led_net_0, 
        sb_sb_0_STAMP_PSELx, MISO_c, MMUART_0_RXD_F2M_c, 
        RXSM_LO_c, RXSM_SODS_c, RXSM_SOE_c, stamp0_ready_dms1_c, 
        stamp0_ready_dms2_c, stamp0_ready_temp_c, 
        stamp0_spi_miso_c, ENABLE_MEMORY_LED_c, LED_HEARTBEAT_c, 
        LED_RECORDING_c, MMUART_0_TXD_M2F_c, MOSI_c, SCLK_c, 
        adc_start_c, nCS1_c, nCS2_c, stamp0_spi_clock_c, 
        stamp0_spi_dms1_cs_c, stamp0_spi_dms2_cs_c, 
        stamp0_spi_temp_cs_c, mosi_cl, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[31]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[30]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[29]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[28]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[27]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[26]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[25]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[24]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[23]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[22]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[21]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[20]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[19]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[18]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[17]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[16]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1]\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0]\, 
        \sb_sb_0/STAMP_PADDRS[15]\, \sb_sb_0/STAMP_PADDRS[14]\, 
        \sb_sb_0/STAMP_PADDRS[13]\, \sb_sb_0/STAMP_PADDRS[12]\, 
        \sb_sb_0/Memory_0_intr_or_0_Y\, 
        \sb_sb_0/FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC\, 
        \sb_sb_0/FIC_0_LOCK\, \sb_sb_0/PREADY_0_iv_i\, 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx\, 
        \sb_sb_0/CoreAPB3_0/iPSELS_raw_1_0_Z[0]\, 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS_Z[2]\, 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS[1]\, 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS[0]\, 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, 
        \sb_sb_0/CCC_0/GL0_net\, \sb_sb_0/CCC_0/GL1_net\, 
        \STAMP_0/component_state_Z[5]\, 
        \STAMP_0/component_state_Z[4]\, 
        \STAMP_0/component_state_Z[3]\, 
        \STAMP_0/component_state_Z[2]\, 
        \STAMP_0/component_state_Z[1]\, 
        \STAMP_0/component_state_Z[0]\, 
        \STAMP_0/async_prescaler_count_Z[11]\, 
        \STAMP_0/async_prescaler_count_Z[10]\, 
        \STAMP_0/async_prescaler_count_Z[9]\, 
        \STAMP_0/async_prescaler_count_Z[8]\, 
        \STAMP_0/async_prescaler_count_Z[7]\, 
        \STAMP_0/async_prescaler_count_Z[6]\, 
        \STAMP_0/async_prescaler_count_Z[5]\, 
        \STAMP_0/async_prescaler_count_Z[4]\, 
        \STAMP_0/async_prescaler_count_Z[3]\, 
        \STAMP_0/async_prescaler_count_Z[2]\, 
        \STAMP_0/async_prescaler_count_Z[1]\, 
        \STAMP_0/async_prescaler_count_Z[0]\, 
        \STAMP_0/async_prescaler_count_5_Z[11]\, 
        \STAMP_0/async_prescaler_count_5_Z[8]\, 
        \STAMP_0/async_prescaler_count_5_Z[7]\, 
        \STAMP_0/async_prescaler_count_5_Z[6]\, 
        \STAMP_0/async_prescaler_count_5_Z[2]\, 
        \STAMP_0/async_prescaler_count_5_Z[0]\, 
        \STAMP_0/spi_rx_data[15]\, \STAMP_0/spi_rx_data[14]\, 
        \STAMP_0/spi_rx_data[13]\, \STAMP_0/spi_rx_data[12]\, 
        \STAMP_0/spi_rx_data[11]\, \STAMP_0/spi_rx_data[10]\, 
        \STAMP_0/spi_rx_data[9]\, \STAMP_0/spi_rx_data[8]\, 
        \STAMP_0/spi_rx_data[7]\, \STAMP_0/spi_rx_data[6]\, 
        \STAMP_0/spi_rx_data[5]\, \STAMP_0/spi_rx_data[4]\, 
        \STAMP_0/spi_rx_data[3]\, \STAMP_0/spi_rx_data[2]\, 
        \STAMP_0/spi_rx_data[1]\, \STAMP_0/spi_rx_data[0]\, 
        \STAMP_0/spi_request_for_Z[1]\, 
        \STAMP_0/spi_request_for_Z[0]\, 
        \STAMP_0/async_state_Z[1]\, \STAMP_0/async_state_Z[0]\, 
        \STAMP_0/async_state_17[1]\, 
        \STAMP_0/un1_spi_rx_data_Z[15]\, 
        \STAMP_0/un1_spi_rx_data_Z[14]\, 
        \STAMP_0/un1_spi_rx_data_Z[13]\, 
        \STAMP_0/un1_spi_rx_data_Z[12]\, 
        \STAMP_0/un1_spi_rx_data_Z[11]\, 
        \STAMP_0/un1_spi_rx_data_Z[10]\, 
        \STAMP_0/un1_spi_rx_data_Z[9]\, 
        \STAMP_0/un1_spi_rx_data_Z[8]\, 
        \STAMP_0/un1_spi_rx_data_Z[7]\, 
        \STAMP_0/un1_spi_rx_data_Z[6]\, 
        \STAMP_0/un1_spi_rx_data_Z[5]\, 
        \STAMP_0/un1_spi_rx_data_Z[4]\, 
        \STAMP_0/un1_spi_rx_data_Z[3]\, 
        \STAMP_0/un1_spi_rx_data_Z[2]\, 
        \STAMP_0/un1_spi_rx_data_Z[1]\, 
        \STAMP_0/un1_spi_rx_data_Z[0]\, \STAMP_0/config_Z[31]\, 
        \STAMP_0/config_Z[30]\, \STAMP_0/config_Z[29]\, 
        \STAMP_0/config_Z[28]\, \STAMP_0/config_Z[27]\, 
        \STAMP_0/config_Z[26]\, \STAMP_0/config_Z[25]\, 
        \STAMP_0/config_Z[24]\, \STAMP_0/config_Z[23]\, 
        \STAMP_0/config_Z[22]\, \STAMP_0/config_Z[21]\, 
        \STAMP_0/config_Z[20]\, \STAMP_0/config_Z[19]\, 
        \STAMP_0/config_Z[18]\, \STAMP_0/config_Z[17]\, 
        \STAMP_0/config_Z[16]\, \STAMP_0/config_Z[15]\, 
        \STAMP_0/config_Z[14]\, \STAMP_0/config_Z[13]\, 
        \STAMP_0/config_Z[12]\, \STAMP_0/config_Z[11]\, 
        \STAMP_0/config_Z[10]\, \STAMP_0/config_Z[9]\, 
        \STAMP_0/config_Z[8]\, \STAMP_0/config_Z[7]\, 
        \STAMP_0/config_Z[6]\, \STAMP_0/config_Z[5]\, 
        \STAMP_0/config_Z[4]\, \STAMP_0/config_Z[3]\, 
        \STAMP_0/config_8[31]\, \STAMP_0/spi_tx_data_Z[15]\, 
        \STAMP_0/spi_tx_data_Z[14]\, \STAMP_0/spi_tx_data_Z[13]\, 
        \STAMP_0/spi_tx_data_Z[12]\, \STAMP_0/spi_tx_data_Z[11]\, 
        \STAMP_0/spi_tx_data_Z[10]\, \STAMP_0/spi_tx_data_Z[9]\, 
        \STAMP_0/spi_tx_data_Z[8]\, \STAMP_0/spi_tx_data_Z[7]\, 
        \STAMP_0/spi_tx_data_Z[6]\, \STAMP_0/spi_tx_data_Z[5]\, 
        \STAMP_0/spi_tx_data_Z[4]\, \STAMP_0/spi_tx_data_Z[3]\, 
        \STAMP_0/spi_tx_data_Z[2]\, \STAMP_0/spi_tx_data_Z[1]\, 
        \STAMP_0/spi_tx_data_Z[0]\, \STAMP_0/un1_pwdata_Z[12]\, 
        \STAMP_0/un1_pwdata_Z[11]\, \STAMP_0/un1_pwdata_Z[10]\, 
        \STAMP_0/dummy_Z[31]\, \STAMP_0/dummy_Z[30]\, 
        \STAMP_0/dummy_Z[29]\, \STAMP_0/dummy_Z[28]\, 
        \STAMP_0/dummy_Z[27]\, \STAMP_0/dummy_Z[26]\, 
        \STAMP_0/dummy_Z[25]\, \STAMP_0/dummy_Z[24]\, 
        \STAMP_0/dummy_Z[23]\, \STAMP_0/dummy_Z[22]\, 
        \STAMP_0/dummy_Z[21]\, \STAMP_0/dummy_Z[20]\, 
        \STAMP_0/dummy_Z[19]\, \STAMP_0/dummy_Z[18]\, 
        \STAMP_0/dummy_Z[17]\, \STAMP_0/dummy_Z[16]\, 
        \STAMP_0/dummy_Z[15]\, \STAMP_0/dummy_Z[14]\, 
        \STAMP_0/dummy_Z[13]\, \STAMP_0/dummy_Z[12]\, 
        \STAMP_0/dummy_Z[11]\, \STAMP_0/dummy_Z[10]\, 
        \STAMP_0/dummy_Z[9]\, \STAMP_0/dummy_Z[8]\, 
        \STAMP_0/dummy_Z[7]\, \STAMP_0/dummy_Z[6]\, 
        \STAMP_0/dummy_Z[5]\, \STAMP_0/dummy_Z[4]\, 
        \STAMP_0/dummy_Z[3]\, \STAMP_0/dummy_Z[2]\, 
        \STAMP_0/dummy_Z[1]\, \STAMP_0/dummy_Z[0]\, 
        \STAMP_0/component_state_ns[3]\, 
        \STAMP_0/component_state_ns[2]\, 
        \STAMP_0/component_state_ns[1]\, 
        \STAMP_0/delay_counter_Z[27]\, 
        \STAMP_0/delay_counter_Z[26]\, 
        \STAMP_0/delay_counter_Z[25]\, 
        \STAMP_0/delay_counter_Z[24]\, 
        \STAMP_0/delay_counter_Z[23]\, 
        \STAMP_0/delay_counter_Z[22]\, 
        \STAMP_0/delay_counter_Z[21]\, 
        \STAMP_0/delay_counter_Z[20]\, 
        \STAMP_0/delay_counter_Z[19]\, 
        \STAMP_0/delay_counter_Z[18]\, 
        \STAMP_0/delay_counter_Z[17]\, 
        \STAMP_0/delay_counter_Z[16]\, 
        \STAMP_0/delay_counter_Z[15]\, 
        \STAMP_0/delay_counter_Z[14]\, 
        \STAMP_0/delay_counter_Z[13]\, 
        \STAMP_0/delay_counter_Z[12]\, 
        \STAMP_0/delay_counter_Z[11]\, 
        \STAMP_0/delay_counter_Z[10]\, 
        \STAMP_0/delay_counter_Z[9]\, 
        \STAMP_0/delay_counter_Z[8]\, 
        \STAMP_0/delay_counter_Z[7]\, 
        \STAMP_0/delay_counter_Z[6]\, 
        \STAMP_0/delay_counter_Z[5]\, 
        \STAMP_0/delay_counter_Z[4]\, 
        \STAMP_0/delay_counter_Z[3]\, 
        \STAMP_0/delay_counter_Z[2]\, 
        \STAMP_0/delay_counter_Z[1]\, 
        \STAMP_0/delay_counter_Z[0]\, 
        \STAMP_0/delay_counter_lm[27]\, 
        \STAMP_0/delay_counter_lm[26]\, 
        \STAMP_0/delay_counter_lm[25]\, 
        \STAMP_0/delay_counter_lm[24]\, 
        \STAMP_0/delay_counter_lm[23]\, 
        \STAMP_0/delay_counter_lm[22]\, 
        \STAMP_0/delay_counter_lm[21]\, 
        \STAMP_0/delay_counter_lm[20]\, 
        \STAMP_0/delay_counter_lm[19]\, 
        \STAMP_0/delay_counter_lm[18]\, 
        \STAMP_0/delay_counter_lm[17]\, 
        \STAMP_0/delay_counter_lm[16]\, 
        \STAMP_0/delay_counter_lm[15]\, 
        \STAMP_0/delay_counter_lm[14]\, 
        \STAMP_0/delay_counter_lm[13]\, 
        \STAMP_0/delay_counter_lm[12]\, 
        \STAMP_0/delay_counter_lm[11]\, 
        \STAMP_0/delay_counter_lm[10]\, 
        \STAMP_0/delay_counter_lm[9]\, 
        \STAMP_0/delay_counter_lm[8]\, 
        \STAMP_0/delay_counter_lm[7]\, 
        \STAMP_0/delay_counter_lm[6]\, 
        \STAMP_0/delay_counter_lm[5]\, 
        \STAMP_0/delay_counter_lm[4]\, 
        \STAMP_0/delay_counter_lm[3]\, 
        \STAMP_0/delay_counter_lm[2]\, 
        \STAMP_0/delay_counter_lm[1]\, 
        \STAMP_0/delay_counter_lm[0]\, 
        \STAMP_0/status_async_cycles_lm[5]\, 
        \STAMP_0/status_async_cycles_lm[4]\, 
        \STAMP_0/status_async_cycles_lm[3]\, 
        \STAMP_0/status_async_cycles_lm[2]\, 
        \STAMP_0/status_async_cycles_lm[1]\, 
        \STAMP_0/status_async_cycles_lm[0]\, 
        \STAMP_0/delay_counter_cry_Z[26]\, 
        \STAMP_0/delay_counter_cry_Z[25]\, 
        \STAMP_0/delay_counter_cry_Z[24]\, 
        \STAMP_0/delay_counter_cry_Z[23]\, 
        \STAMP_0/delay_counter_cry_Z[22]\, 
        \STAMP_0/delay_counter_cry_Z[21]\, 
        \STAMP_0/delay_counter_cry_Z[20]\, 
        \STAMP_0/delay_counter_cry_Z[19]\, 
        \STAMP_0/delay_counter_cry_Z[18]\, 
        \STAMP_0/delay_counter_cry_Z[17]\, 
        \STAMP_0/delay_counter_cry_Z[16]\, 
        \STAMP_0/delay_counter_cry_Z[15]\, 
        \STAMP_0/delay_counter_cry_Z[14]\, 
        \STAMP_0/delay_counter_cry_Z[13]\, 
        \STAMP_0/delay_counter_cry_Z[12]\, 
        \STAMP_0/delay_counter_cry_Z[11]\, 
        \STAMP_0/delay_counter_cry_Z[10]\, 
        \STAMP_0/delay_counter_cry_Z[9]\, 
        \STAMP_0/delay_counter_cry_Z[8]\, 
        \STAMP_0/delay_counter_cry_Z[7]\, 
        \STAMP_0/delay_counter_cry_Z[6]\, 
        \STAMP_0/delay_counter_cry_Z[5]\, 
        \STAMP_0/delay_counter_cry_Z[4]\, 
        \STAMP_0/delay_counter_cry_Z[3]\, 
        \STAMP_0/delay_counter_cry_Z[2]\, 
        \STAMP_0/delay_counter_cry_Z[1]\, 
        \STAMP_0/delay_counter_cry_Z[0]\, 
        \STAMP_0/delay_counter_cry_Y[0]\, 
        \STAMP_0/delay_counter_s[26]\, 
        \STAMP_0/delay_counter_s[25]\, 
        \STAMP_0/delay_counter_s[24]\, 
        \STAMP_0/delay_counter_s[23]\, 
        \STAMP_0/delay_counter_s[22]\, 
        \STAMP_0/delay_counter_s[21]\, 
        \STAMP_0/delay_counter_s[20]\, 
        \STAMP_0/delay_counter_s[19]\, 
        \STAMP_0/delay_counter_s[18]\, 
        \STAMP_0/delay_counter_s[17]\, 
        \STAMP_0/delay_counter_s[16]\, 
        \STAMP_0/delay_counter_s[15]\, 
        \STAMP_0/delay_counter_s[14]\, 
        \STAMP_0/delay_counter_s[13]\, 
        \STAMP_0/delay_counter_s[12]\, 
        \STAMP_0/delay_counter_s[11]\, 
        \STAMP_0/delay_counter_s[10]\, 
        \STAMP_0/delay_counter_s[9]\, 
        \STAMP_0/delay_counter_s[8]\, 
        \STAMP_0/delay_counter_s[7]\, 
        \STAMP_0/delay_counter_s[6]\, 
        \STAMP_0/delay_counter_s[5]\, 
        \STAMP_0/delay_counter_s[4]\, 
        \STAMP_0/delay_counter_s[3]\, 
        \STAMP_0/delay_counter_s[2]\, 
        \STAMP_0/delay_counter_s[1]\, 
        \STAMP_0/delay_counter_s_Z[27]\, 
        \STAMP_0/status_async_cycles_cry_Z[4]\, 
        \STAMP_0/status_async_cycles_cry_Z[3]\, 
        \STAMP_0/status_async_cycles_cry_Z[2]\, 
        \STAMP_0/status_async_cycles_cry_Z[1]\, 
        \STAMP_0/status_async_cycles_s[4]\, 
        \STAMP_0/status_async_cycles_s[3]\, 
        \STAMP_0/status_async_cycles_s[2]\, 
        \STAMP_0/status_async_cycles_s[1]\, 
        \STAMP_0/status_async_cycles_s_Z[5]\, 
        \STAMP_0/un1_spi_rx_data_2_1_0_Z[2]\, 
        \STAMP_0/un1_spi_rx_data_2_1_0_Z[1]\, 
        \STAMP_0/un1_spi_rx_data_2_1_0_Z[0]\, 
        \STAMP_0/component_state_ns_0_1_Z[3]\, 
        \STAMP_0/component_state_ns_0_0_a3_1_Z[2]\, 
        \STAMP_0/component_state_ns_0_0_0_Z[2]\, 
        \STAMP_0/component_state_ns_0_0_0_Z[1]\, 
        \STAMP_0/component_state_ns_0_i_0_tz_Z[0]\, 
        \STAMP_0/component_state_RNIFR114_Z[0]\, 
        \STAMP_0/component_state_ns_0_i_a3_1_1_Z[0]\, 
        \STAMP_0/component_state_ns_0_i_0_0_Z[0]\, 
        \STAMP_0/stamp0_ready_temp_c_i\, 
        \STAMP_0/stamp0_ready_dms2_c_i\, 
        \STAMP_0/stamp0_ready_dms1_c_i\, 
        \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, 
        \STAMP_0/un5_async_prescaler_count_cry_4_S\, 
        \STAMP_0/un5_async_prescaler_count_cry_5_S\, 
        \STAMP_0/un5_async_prescaler_count_cry_9_S\, 
        \STAMP_0/un5_async_prescaler_count_cry_10_S\, 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, \STAMP_0/N_567_i\, 
        \STAMP_0/un1_presetn_inv_4_i_0_Z\, \STAMP_0/N_568_i\, 
        \STAMP_0/N_90_i\, 
        \STAMP_0/un5_async_prescaler_count_cry_1_S\, 
        \STAMP_0/un5_async_prescaler_count_cry_3_S\, 
        \STAMP_0/measurement_dms2_1_sqmuxa\, 
        \STAMP_0/measurement_temp_1_sqmuxa\, \STAMP_0/N_119_i\, 
        \STAMP_0/un1_presetn_inv_i\, \STAMP_0/config_143\, 
        \STAMP_0/un1_component_state_6_i\, \STAMP_0/N_297_i\, 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, \STAMP_0/N_296_i\, 
        \STAMP_0/N_295_i\, \STAMP_0/N_294_i\, \STAMP_0/N_293_i\, 
        \STAMP_0/N_292_i\, \STAMP_0/N_291_i\, \STAMP_0/N_290_i\, 
        \STAMP_0/N_289_i\, \STAMP_0/N_266_i\, \STAMP_0/N_267_i\, 
        \STAMP_0/N_268_i\, 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, 
        \STAMP_0/N_298_i\, \STAMP_0/N_116_i\, 
        \STAMP_0/un1_drdy_flank_detected_dms1_0_sqmuxa_1_Z\, 
        \STAMP_0/drdy_flank_detected_dms1_0_sqmuxa_1\, 
        \STAMP_0/apb_is_reset_Z\, 
        \STAMP_0/apb_is_atomic_0_sqmuxa\, 
        \STAMP_0/apb_is_atomic_Z\, 
        \STAMP_0/spi_dms2_cs_13_iv_i_Z\, \STAMP_0/N_46\, 
        \STAMP_0/spi_temp_cs_13_iv_i_Z\, 
        \STAMP_0/un1_component_state_13_i_0_Z\, 
        \STAMP_0/spi_dms1_cs_14_iv_i_Z\, 
        \STAMP_0/un1_component_state_14_i_0_Z\, 
        \STAMP_0/apb_spi_finished_Z\, 
        \STAMP_0/un1_apb_spi_finished_1_f0_Z\, 
        \STAMP_0/PREADY_0_sqmuxa_2\, 
        \STAMP_0/un1_PREADY_0_sqmuxa_3_0_Z\, 
        \STAMP_0/drdy_flank_detected_temp_Z\, 
        \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_2_i_Z\, 
        \STAMP_0/drdy_flank_detected_dms2_Z\, 
        \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_2_i_Z\, 
        \STAMP_0/drdy_flank_detected_dms1_Z\, 
        \STAMP_0/drdy_flank_detected_dms1_1_sqmuxa_1_i_Z\, 
        \STAMP_0/enable\, \STAMP_0/spi_enable_RNO_Z\, 
        \STAMP_0/N_244\, \STAMP_0/new_avail_0_sqmuxa_1\, 
        \STAMP_0/un1_new_avail_1_sqmuxa_3_i_0_Z\, 
        \STAMP_0/request_resync_1_sqmuxa_1_Z\, \STAMP_0/N_152\, 
        \STAMP_0/status_temp_overwrittenVal_9_Z\, 
        \STAMP_0/un1_new_avail_0_sqmuxa_2_Z\, 
        \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_1\, 
        \STAMP_0/N_117_i\, \STAMP_0/un1_new_avail_0_sqmuxa_3_Z\, 
        \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_1\, 
        \STAMP_0/N_100_i\, \STAMP_0/N_536_i\, \STAMP_0/N_487_i\, 
        \STAMP_0/N_678\, \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, 
        \STAMP_0/N_679\, \STAMP_0/N_681\, \STAMP_0/N_666\, 
        \STAMP_0/N_667\, \STAMP_0/N_668\, \STAMP_0/N_669\, 
        \STAMP_0/N_670\, \STAMP_0/N_671\, \STAMP_0/N_672\, 
        \STAMP_0/N_673\, \STAMP_0/N_674\, \STAMP_0/N_675\, 
        \STAMP_0/N_676\, \STAMP_0/N_677\, \STAMP_0/N_118_i\, 
        \STAMP_0/status_async_cycles_1_sqmuxa_1_i_Z\, 
        \STAMP_0/un45_async_state_cry_0_Z\, 
        \STAMP_0/un45_async_state_cry_1_Z\, 
        \STAMP_0/un45_async_state_cry_2_Z\, 
        \STAMP_0/un45_async_state_cry_3_Z\, 
        \STAMP_0/un45_async_state_cry_4_Z\, 
        \STAMP_0/un45_async_state_cry_5_Z\, 
        \STAMP_0/status_async_cycles_s_388_FCO\, 
        \STAMP_0/un5_async_prescaler_count_s_1_391_FCO\, 
        \STAMP_0/un5_async_prescaler_count_cry_1_Z\, 
        \STAMP_0/un5_async_prescaler_count_cry_2_Z\, 
        \STAMP_0/un5_async_prescaler_count_cry_2_S\, 
        \STAMP_0/un5_async_prescaler_count_cry_3_Z\, 
        \STAMP_0/un5_async_prescaler_count_cry_4_Z\, 
        \STAMP_0/un5_async_prescaler_count_cry_5_Z\, 
        \STAMP_0/un5_async_prescaler_count_cry_6_Z\, 
        \STAMP_0/un5_async_prescaler_count_cry_6_S\, 
        \STAMP_0/un5_async_prescaler_count_cry_7_Z\, 
        \STAMP_0/un5_async_prescaler_count_cry_7_S\, 
        \STAMP_0/un5_async_prescaler_count_cry_8_Z\, 
        \STAMP_0/un5_async_prescaler_count_cry_8_S\, 
        \STAMP_0/un5_async_prescaler_count_cry_9_Z\, 
        \STAMP_0/un5_async_prescaler_count_s_11_S\, 
        \STAMP_0/un5_async_prescaler_count_cry_10_Z\, 
        \STAMP_0/N_109_i\, \STAMP_0/N_329\, 
        \STAMP_0/un1_new_avail_0_sqmuxa_1\, \STAMP_0/N_160\, 
        \STAMP_0/N_168\, \STAMP_0/N_650\, \STAMP_0/N_651\, 
        \STAMP_0/N_652\, \STAMP_0/un27_paddr_i_0\, 
        \STAMP_0/un13_paddr_i_0\, 
        \STAMP_0/un1_spi_rx_data_sn_N_5\, 
        \STAMP_0/apb_spi_finished_0_sqmuxa\, \STAMP_0/N_158\, 
        \STAMP_0/spi_busy\, \STAMP_0/N_111_i\, \STAMP_0/N_164\, 
        \STAMP_0/N_110_i\, \STAMP_0/N_165\, \STAMP_0/N_112_i\, 
        \STAMP_0/N_166\, \STAMP_0/request_resync_0_sqmuxa\, 
        \STAMP_0/un52_paddr_5_Z\, \STAMP_0/un52_paddr_2_Z\, 
        \STAMP_0/N_596\, \STAMP_0/N_614\, \STAMP_0/N_611\, 
        \STAMP_0/N_589\, \STAMP_0/N_587\, \STAMP_0/N_610\, 
        \STAMP_0/N_609\, \STAMP_0/N_608\, \STAMP_0/N_607\, 
        \STAMP_0/N_606\, \STAMP_0/N_605\, \STAMP_0/N_604\, 
        \STAMP_0/N_603\, \STAMP_0/N_602\, \STAMP_0/N_601\, 
        \STAMP_0/N_600\, \STAMP_0/N_599\, \STAMP_0/N_598\, 
        \STAMP_0/N_597\, \STAMP_0/N_595\, \STAMP_0/N_594\, 
        \STAMP_0/N_593\, \STAMP_0/N_592\, \STAMP_0/N_591\, 
        \STAMP_0/N_590\, \STAMP_0/N_588\, \STAMP_0/N_586\, 
        \STAMP_0/N_218\, \STAMP_0/N_612\, 
        \STAMP_0/un1_component_state_8_0_Z\, 
        \STAMP_0/dummy_1_sqmuxa_2_Z\, \STAMP_0/un60_paddr_3_2_Z\, 
        \STAMP_0/un27_paddr_1_Z\, 
        \STAMP_0/async_state_0_sqmuxa_1_1_Z\, 
        \STAMP_0/N_517_i_0_a2_20\, \STAMP_0/N_517_i_0_a2_19\, 
        \STAMP_0/N_517_i_0_a2_18\, \STAMP_0/N_517_i_0_a2_17\, 
        \STAMP_0/N_517_i_0_a2_16\, \STAMP_0/N_517_i_0_a2_15\, 
        \STAMP_0/N_517_i_0_a2_14\, 
        \STAMP_0/un1_async_prescaler_countlt8\, 
        \STAMP_0/un52_paddr_2_0_Z\, 
        \STAMP_0/apb_spi_finished_1_sqmuxa\, 
        \STAMP_0/apb_spi_finished_0_sqmuxa_1\, \STAMP_0/N_162_i\, 
        \STAMP_0/N_155\, \STAMP_0/N_156\, \STAMP_0/N_163\, 
        \STAMP_0/N_167\, \STAMP_0/N_219\, 
        \STAMP_0/async_state_0_sqmuxa_Z\, 
        \STAMP_0/spi_request_for_2_sqmuxa\, 
        \STAMP_0/spi_dms2_cs_1_sqmuxa_1\, \STAMP_0/N_216_i\, 
        \STAMP_0/N_620\, \STAMP_0/N_626\, \STAMP_0/N_627\, 
        \STAMP_0/N_628\, \STAMP_0/N_629\, \STAMP_0/N_631\, 
        \STAMP_0/N_632\, \STAMP_0/N_633\, \STAMP_0/N_634\, 
        \STAMP_0/N_635\, \STAMP_0/N_636\, \STAMP_0/N_637\, 
        \STAMP_0/N_638\, \STAMP_0/N_639\, \STAMP_0/N_640\, 
        \STAMP_0/N_641\, \STAMP_0/N_642\, \STAMP_0/N_643\, 
        \STAMP_0/N_644\, \STAMP_0/N_630\, 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, \STAMP_0/N_648\, 
        \STAMP_0/N_645\, \STAMP_0/N_623\, \STAMP_0/N_621\, 
        \STAMP_0/N_625\, \STAMP_0/N_624\, \STAMP_0/N_622\, 
        \STAMP_0/N_220\, \STAMP_0/N_646\, 
        \STAMP_0/un1_component_state_9_i_a3_1_Z\, 
        \STAMP_0/un76_paddr_0_a2_2_Z\, \STAMP_0/un52_paddr_2_1\, 
        \STAMP_0/dummy_1_sqmuxa_4_Z\, 
        \STAMP_0/un1_async_prescaler_countlt10\, 
        \STAMP_0/un68_paddr_1_0_Z\, 
        \STAMP_0/spi_dms1_cs_0_sqmuxa_3\, 
        \STAMP_0/N_517_i_0_a2_25\, \STAMP_0/N_337\, 
        \STAMP_0/un1_async_state_0_sqmuxa_i\, 
        \STAMP_0/un76_paddr\, \STAMP_0/un85_paddr_3_0_tz_Z\, 
        \STAMP_0/N_663\, \STAMP_0/N_656\, \STAMP_0/N_654\, 
        \STAMP_0/N_665\, \STAMP_0/N_664\, \STAMP_0/N_662\, 
        \STAMP_0/N_661\, \STAMP_0/N_660\, \STAMP_0/N_659\, 
        \STAMP_0/N_658\, \STAMP_0/N_657\, \STAMP_0/N_655\, 
        \STAMP_0/N_653\, \STAMP_0/N_238\, \STAMP_0/N_364\, 
        \STAMP_0/un1_async_prescaler_count\, 
        \STAMP_0/un85_paddr_3_Z\, \STAMP_0/N_353\, 
        \STAMP_0/N_263\, \STAMP_0/N_331\, \STAMP_0/N_333\, 
        \STAMP_0/N_363\, \STAMP_0/status_async_cycles_1_sqmuxa_Z\, 
        \STAMP_0/un1_component_state_13_i_a3_0_0_Z\, 
        \STAMP_0/un1_presetn_inv_Z\, \STAMP_0/N_215\, 
        \STAMP_0/status_async_cycles_3_sqmuxa\, 
        \STAMP_0/status_async_cycles_2_sqmuxa\, \STAMP_0/N_361\, 
        \STAMP_0/N_248_2\, \STAMP_0/N_197\, \STAMP_0/N_204\, 
        \STAMP_0/N_206\, \STAMP_0/spi/rx_buffer_Z[15]\, 
        \STAMP_0/spi/rx_buffer_Z[14]\, 
        \STAMP_0/spi/rx_buffer_Z[13]\, 
        \STAMP_0/spi/rx_buffer_Z[12]\, 
        \STAMP_0/spi/rx_buffer_Z[11]\, 
        \STAMP_0/spi/rx_buffer_Z[10]\, 
        \STAMP_0/spi/rx_buffer_Z[9]\, 
        \STAMP_0/spi/rx_buffer_Z[8]\, 
        \STAMP_0/spi/rx_buffer_Z[7]\, 
        \STAMP_0/spi/rx_buffer_Z[6]\, 
        \STAMP_0/spi/rx_buffer_Z[5]\, 
        \STAMP_0/spi/rx_buffer_Z[4]\, 
        \STAMP_0/spi/rx_buffer_Z[3]\, 
        \STAMP_0/spi/rx_buffer_Z[2]\, 
        \STAMP_0/spi/rx_buffer_Z[1]\, 
        \STAMP_0/spi/rx_buffer_Z[0]\, 
        \STAMP_0/spi/tx_buffer_Z[15]\, 
        \STAMP_0/spi/tx_buffer_Z[14]\, 
        \STAMP_0/spi/tx_buffer_Z[13]\, 
        \STAMP_0/spi/tx_buffer_Z[12]\, 
        \STAMP_0/spi/tx_buffer_Z[11]\, 
        \STAMP_0/spi/tx_buffer_Z[10]\, 
        \STAMP_0/spi/tx_buffer_Z[9]\, 
        \STAMP_0/spi/tx_buffer_Z[8]\, 
        \STAMP_0/spi/tx_buffer_Z[7]\, 
        \STAMP_0/spi/tx_buffer_Z[6]\, 
        \STAMP_0/spi/tx_buffer_Z[5]\, 
        \STAMP_0/spi/tx_buffer_Z[4]\, 
        \STAMP_0/spi/tx_buffer_Z[3]\, 
        \STAMP_0/spi/tx_buffer_Z[2]\, 
        \STAMP_0/spi/tx_buffer_Z[1]\, 
        \STAMP_0/spi/tx_buffer_Z[0]\, 
        \STAMP_0/spi/ss_n_buffer_Z[0]\, \STAMP_0/spi/state_Z[0]\, 
        \STAMP_0/spi/clk_toggles_Z[5]\, 
        \STAMP_0/spi/clk_toggles_Z[4]\, 
        \STAMP_0/spi/clk_toggles_Z[3]\, 
        \STAMP_0/spi/clk_toggles_Z[2]\, 
        \STAMP_0/spi/clk_toggles_Z[1]\, 
        \STAMP_0/spi/clk_toggles_Z[0]\, 
        \STAMP_0/spi/clk_toggles_lm[5]\, 
        \STAMP_0/spi/clk_toggles_lm[4]\, 
        \STAMP_0/spi/clk_toggles_lm[3]\, 
        \STAMP_0/spi/clk_toggles_lm[2]\, 
        \STAMP_0/spi/clk_toggles_lm[1]\, 
        \STAMP_0/spi/clk_toggles_lm[0]\, 
        \STAMP_0/spi/count_Z[31]\, \STAMP_0/spi/count_Z[30]\, 
        \STAMP_0/spi/count_Z[29]\, \STAMP_0/spi/count_Z[28]\, 
        \STAMP_0/spi/count_Z[27]\, \STAMP_0/spi/count_Z[26]\, 
        \STAMP_0/spi/count_Z[25]\, \STAMP_0/spi/count_Z[24]\, 
        \STAMP_0/spi/count_Z[23]\, \STAMP_0/spi/count_Z[22]\, 
        \STAMP_0/spi/count_Z[21]\, \STAMP_0/spi/count_Z[20]\, 
        \STAMP_0/spi/count_Z[19]\, \STAMP_0/spi/count_Z[18]\, 
        \STAMP_0/spi/count_Z[17]\, \STAMP_0/spi/count_Z[16]\, 
        \STAMP_0/spi/count_Z[15]\, \STAMP_0/spi/count_Z[14]\, 
        \STAMP_0/spi/count_Z[13]\, \STAMP_0/spi/count_Z[12]\, 
        \STAMP_0/spi/count_Z[11]\, \STAMP_0/spi/count_Z[10]\, 
        \STAMP_0/spi/count_Z[9]\, \STAMP_0/spi/count_Z[8]\, 
        \STAMP_0/spi/count_Z[7]\, \STAMP_0/spi/count_Z[6]\, 
        \STAMP_0/spi/count_Z[5]\, \STAMP_0/spi/count_Z[4]\, 
        \STAMP_0/spi/count_Z[3]\, \STAMP_0/spi/count_Z[2]\, 
        \STAMP_0/spi/count_Z[1]\, \STAMP_0/spi/count_Z[0]\, 
        \STAMP_0/spi/count_lm[31]\, \STAMP_0/spi/count_lm[30]\, 
        \STAMP_0/spi/count_lm[29]\, \STAMP_0/spi/count_lm[28]\, 
        \STAMP_0/spi/count_lm[27]\, \STAMP_0/spi/count_lm[26]\, 
        \STAMP_0/spi/count_lm[25]\, \STAMP_0/spi/count_lm[24]\, 
        \STAMP_0/spi/count_lm[23]\, \STAMP_0/spi/count_lm[22]\, 
        \STAMP_0/spi/count_lm[21]\, \STAMP_0/spi/count_lm[20]\, 
        \STAMP_0/spi/count_lm[19]\, \STAMP_0/spi/count_lm[18]\, 
        \STAMP_0/spi/count_lm[17]\, \STAMP_0/spi/count_lm[16]\, 
        \STAMP_0/spi/count_lm[15]\, \STAMP_0/spi/count_lm[14]\, 
        \STAMP_0/spi/count_lm[13]\, \STAMP_0/spi/count_lm[12]\, 
        \STAMP_0/spi/count_lm[11]\, \STAMP_0/spi/count_lm[10]\, 
        \STAMP_0/spi/count_lm[9]\, \STAMP_0/spi/count_lm[8]\, 
        \STAMP_0/spi/count_lm[7]\, \STAMP_0/spi/count_lm[6]\, 
        \STAMP_0/spi/count_lm[5]\, \STAMP_0/spi/count_lm[4]\, 
        \STAMP_0/spi/count_lm[3]\, \STAMP_0/spi/count_lm[2]\, 
        \STAMP_0/spi/count_lm[1]\, \STAMP_0/spi/count_lm[0]\, 
        \STAMP_0/spi/count_cry_Z[30]\, 
        \STAMP_0/spi/count_cry_Z[29]\, 
        \STAMP_0/spi/count_cry_Z[28]\, 
        \STAMP_0/spi/count_cry_Z[27]\, 
        \STAMP_0/spi/count_cry_Z[26]\, 
        \STAMP_0/spi/count_cry_Z[25]\, 
        \STAMP_0/spi/count_cry_Z[24]\, 
        \STAMP_0/spi/count_cry_Z[23]\, 
        \STAMP_0/spi/count_cry_Z[22]\, 
        \STAMP_0/spi/count_cry_Z[21]\, 
        \STAMP_0/spi/count_cry_Z[20]\, 
        \STAMP_0/spi/count_cry_Z[19]\, 
        \STAMP_0/spi/count_cry_Z[18]\, 
        \STAMP_0/spi/count_cry_Z[17]\, 
        \STAMP_0/spi/count_cry_Z[16]\, 
        \STAMP_0/spi/count_cry_Z[15]\, 
        \STAMP_0/spi/count_cry_Z[14]\, 
        \STAMP_0/spi/count_cry_Z[13]\, 
        \STAMP_0/spi/count_cry_Z[12]\, 
        \STAMP_0/spi/count_cry_Z[11]\, 
        \STAMP_0/spi/count_cry_Z[10]\, 
        \STAMP_0/spi/count_cry_Z[9]\, 
        \STAMP_0/spi/count_cry_Z[8]\, 
        \STAMP_0/spi/count_cry_Z[7]\, 
        \STAMP_0/spi/count_cry_Z[6]\, 
        \STAMP_0/spi/count_cry_Z[5]\, 
        \STAMP_0/spi/count_cry_Z[4]\, 
        \STAMP_0/spi/count_cry_Z[3]\, 
        \STAMP_0/spi/count_cry_Z[2]\, 
        \STAMP_0/spi/count_cry_Z[1]\, \STAMP_0/spi/count_s[30]\, 
        \STAMP_0/spi/count_s[29]\, \STAMP_0/spi/count_s[28]\, 
        \STAMP_0/spi/count_s[27]\, \STAMP_0/spi/count_s[26]\, 
        \STAMP_0/spi/count_s[25]\, \STAMP_0/spi/count_s[24]\, 
        \STAMP_0/spi/count_s[23]\, \STAMP_0/spi/count_s[22]\, 
        \STAMP_0/spi/count_s[21]\, \STAMP_0/spi/count_s[20]\, 
        \STAMP_0/spi/count_s[19]\, \STAMP_0/spi/count_s[18]\, 
        \STAMP_0/spi/count_s[17]\, \STAMP_0/spi/count_s[16]\, 
        \STAMP_0/spi/count_s[15]\, \STAMP_0/spi/count_s[14]\, 
        \STAMP_0/spi/count_s[13]\, \STAMP_0/spi/count_s[12]\, 
        \STAMP_0/spi/count_s[11]\, \STAMP_0/spi/count_s[10]\, 
        \STAMP_0/spi/count_s[9]\, \STAMP_0/spi/count_s[8]\, 
        \STAMP_0/spi/count_s[7]\, \STAMP_0/spi/count_s[6]\, 
        \STAMP_0/spi/count_s[5]\, \STAMP_0/spi/count_s[4]\, 
        \STAMP_0/spi/count_s[3]\, \STAMP_0/spi/count_s[2]\, 
        \STAMP_0/spi/count_s[1]\, \STAMP_0/spi/count_s_Z[31]\, 
        \STAMP_0/spi/clk_toggles_cry_Z[4]\, 
        \STAMP_0/spi/clk_toggles_cry_Z[3]\, 
        \STAMP_0/spi/clk_toggles_cry_Z[2]\, 
        \STAMP_0/spi/clk_toggles_cry_Z[1]\, 
        \STAMP_0/spi/clk_toggles_s[4]\, 
        \STAMP_0/spi/clk_toggles_s[3]\, 
        \STAMP_0/spi/clk_toggles_s[2]\, 
        \STAMP_0/spi/clk_toggles_s[1]\, 
        \STAMP_0/spi/clk_toggles_s_Z[5]\, 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, \STAMP_0/spi/N_140\, 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, \STAMP_0/spi/N_138\, 
        \STAMP_0/spi/N_136\, \STAMP_0/spi/N_134\, 
        \STAMP_0/spi/N_132\, \STAMP_0/spi/N_130\, 
        \STAMP_0/spi/N_128\, \STAMP_0/spi/N_127\, 
        \STAMP_0/spi/N_126\, \STAMP_0/spi/N_125\, 
        \STAMP_0/spi/N_124\, \STAMP_0/spi/N_123\, 
        \STAMP_0/spi/N_122\, \STAMP_0/spi/N_121\, 
        \STAMP_0/spi/N_120\, \STAMP_0/spi/N_50_i\, 
        \STAMP_0/spi/N_333\, \STAMP_0/spi/N_20_i\, 
        \STAMP_0/spi/assert_data_Z\, \STAMP_0/spi/assert_data_5\, 
        \STAMP_0/spi/mosi_1_1\, 
        \STAMP_0/spi/ss_n_buffer_1_sqmuxa\, \STAMP_0/spi/busy_7\, 
        \STAMP_0/spi/N_25_i\, \STAMP_0/spi/N_37_i\, 
        \STAMP_0/spi/N_49_i\, \STAMP_0/spi/count_s_389_FCO\, 
        \STAMP_0/spi/clk_toggles_s_390_FCO\, 
        \STAMP_0/spi/un7_count_NE_i\, 
        \STAMP_0/spi/un7_count_NE_13_Z\, 
        \STAMP_0/spi/un10_count_0_a2_0_0_Z\, 
        \STAMP_0/spi/un10_count_0_a2_0_Z\, 
        \STAMP_0/spi/un7_count_NE_23_Z\, 
        \STAMP_0/spi/un7_count_NE_21_Z\, 
        \STAMP_0/spi/un7_count_NE_20_Z\, 
        \STAMP_0/spi/un7_count_NE_19_Z\, 
        \STAMP_0/spi/un7_count_NE_18_Z\, 
        \STAMP_0/spi/un7_count_NE_17_Z\, 
        \STAMP_0/spi/un7_count_NE_16_Z\, 
        \STAMP_0/spi/un10_count_i\, \STAMP_0/spi/count_0_sqmuxa\, 
        \STAMP_0/spi/N_63\, \STAMP_0/spi/mosi_1_1_2\, 
        \STAMP_0/spi/un7_count_NE_27_Z\, 
        \STAMP_0/spi/un7_count_NE_28_Z\, \STAMP_0/spi/N_30\, 
        \STAMP_0/spi/sclk_buffer_0_sqmuxa\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_i_i_a2_fast_Z[0]\, 
        \MemorySynchronizer_0/temp_1[30]\, 
        \MemorySynchronizer_0/temp_1[29]\, 
        \MemorySynchronizer_0/temp_1[28]\, 
        \MemorySynchronizer_0/temp_1[27]\, 
        \MemorySynchronizer_0/temp_1[26]\, 
        \MemorySynchronizer_0/temp_1[25]\, 
        \MemorySynchronizer_0/temp_1[24]\, 
        \MemorySynchronizer_0/temp_1[23]\, 
        \MemorySynchronizer_0/temp_1[22]\, 
        \MemorySynchronizer_0/temp_1[21]\, 
        \MemorySynchronizer_0/temp_1[20]\, 
        \MemorySynchronizer_0/temp_1[19]\, 
        \MemorySynchronizer_0/temp_1[18]\, 
        \MemorySynchronizer_0/temp_1[17]\, 
        \MemorySynchronizer_0/temp_1[16]\, 
        \MemorySynchronizer_0/temp_1[15]\, 
        \MemorySynchronizer_0/temp_1[14]\, 
        \MemorySynchronizer_0/temp_1[13]\, 
        \MemorySynchronizer_0/temp_1[12]\, 
        \MemorySynchronizer_0/temp_1[11]\, 
        \MemorySynchronizer_0/temp_1[10]\, 
        \MemorySynchronizer_0/temp_1[9]\, 
        \MemorySynchronizer_0/temp_1[8]\, 
        \MemorySynchronizer_0/temp_1[7]\, 
        \MemorySynchronizer_0/temp_1[6]\, 
        \MemorySynchronizer_0/temp_1[5]\, 
        \MemorySynchronizer_0/temp_1[4]\, 
        \MemorySynchronizer_0/temp_1[3]\, 
        \MemorySynchronizer_0/temp_1[2]\, 
        \MemorySynchronizer_0/temp_1[1]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[30]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[29]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[28]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[27]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[26]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[25]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[24]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[23]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[22]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[21]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[19]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[18]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[17]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[16]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[15]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[14]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[13]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[12]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[11]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[10]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[9]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[8]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[7]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[6]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[4]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[3]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[2]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[1]\, 
        \MemorySynchronizer_0/SynchStatusReg2_Z[0]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[30]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[29]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[27]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[25]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[24]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[22]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[19]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[18]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[17]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[15]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[14]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[13]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[12]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[10]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[8]\, 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[7]\, 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[28]\, 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[26]\, 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[23]\, 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[21]\, 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[16]\, 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[11]\, 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[9]\, 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[6]\, 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[2]\, 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[1]\, 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[0]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[31]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[30]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[29]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[28]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[27]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[26]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[25]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[24]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[23]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[22]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[13]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[7]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[6]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[5]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[4]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[3]\, 
        \MemorySynchronizer_0/SynchStatusReg_Z[2]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_34_Z[20]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[30]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[29]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[28]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[27]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[26]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[25]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[24]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[23]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[22]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[21]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[20]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[19]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[18]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[17]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[16]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[15]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[14]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[13]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[12]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[11]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[10]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[9]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[8]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[7]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[6]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[5]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[4]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[3]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[2]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[1]\, 
        \MemorySynchronizer_0/resynctimercounter_Z[0]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[31]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[29]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[27]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[26]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[25]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[24]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[23]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[22]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[21]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[20]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[19]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[18]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[17]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[15]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[14]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[12]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[11]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[10]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[9]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[7]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[5]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[3]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[2]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[0]\, 
        \MemorySynchronizer_0/APBState_Z[1]\, 
        \MemorySynchronizer_0/APBState_Z[0]\, 
        \MemorySynchronizer_0/PRDATA_21[30]\, 
        \MemorySynchronizer_0/PRDATA_21[28]\, 
        \MemorySynchronizer_0/PRDATA_21[16]\, 
        \MemorySynchronizer_0/PRDATA_21[13]\, 
        \MemorySynchronizer_0/PRDATA_21[8]\, 
        \MemorySynchronizer_0/PRDATA_21[6]\, 
        \MemorySynchronizer_0/PRDATA_21[4]\, 
        \MemorySynchronizer_0/PRDATA_21[1]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[31]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[30]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[29]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[28]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[27]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[26]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[25]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[24]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[23]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[22]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[21]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[20]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[19]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[18]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[17]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[16]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[15]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[14]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[13]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[12]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[11]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[10]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[9]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[8]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[7]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[6]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[5]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[4]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[3]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[2]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[1]\, 
        \MemorySynchronizer_0/TimeStampReg_Z[0]\, 
        \MemorySynchronizer_0/TimeStampValue[31]\, 
        \MemorySynchronizer_0/TimeStampValue[30]\, 
        \MemorySynchronizer_0/TimeStampValue[29]\, 
        \MemorySynchronizer_0/TimeStampValue[28]\, 
        \MemorySynchronizer_0/TimeStampValue[27]\, 
        \MemorySynchronizer_0/TimeStampValue[26]\, 
        \MemorySynchronizer_0/TimeStampValue[25]\, 
        \MemorySynchronizer_0/TimeStampValue[24]\, 
        \MemorySynchronizer_0/TimeStampValue[23]\, 
        \MemorySynchronizer_0/TimeStampValue[22]\, 
        \MemorySynchronizer_0/TimeStampValue[21]\, 
        \MemorySynchronizer_0/TimeStampValue[20]\, 
        \MemorySynchronizer_0/TimeStampValue[19]\, 
        \MemorySynchronizer_0/TimeStampValue[18]\, 
        \MemorySynchronizer_0/TimeStampValue[17]\, 
        \MemorySynchronizer_0/TimeStampValue[16]\, 
        \MemorySynchronizer_0/TimeStampValue[15]\, 
        \MemorySynchronizer_0/TimeStampValue[14]\, 
        \MemorySynchronizer_0/TimeStampValue[13]\, 
        \MemorySynchronizer_0/TimeStampValue[12]\, 
        \MemorySynchronizer_0/TimeStampValue[11]\, 
        \MemorySynchronizer_0/TimeStampValue[10]\, 
        \MemorySynchronizer_0/TimeStampValue[9]\, 
        \MemorySynchronizer_0/TimeStampValue[8]\, 
        \MemorySynchronizer_0/TimeStampValue[7]\, 
        \MemorySynchronizer_0/TimeStampValue[6]\, 
        \MemorySynchronizer_0/TimeStampValue[5]\, 
        \MemorySynchronizer_0/TimeStampValue[4]\, 
        \MemorySynchronizer_0/TimeStampValue[3]\, 
        \MemorySynchronizer_0/TimeStampValue[2]\, 
        \MemorySynchronizer_0/TimeStampValue[1]\, 
        \MemorySynchronizer_0/TimeStampValue[0]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        \MemorySynchronizer_0/SynchStatusReg_168[11]\, 
        \MemorySynchronizer_0/SynchStatusReg_168[5]\, 
        \MemorySynchronizer_0/SynchStatusReg_168[4]\, 
        \MemorySynchronizer_0/SynchStatusReg_168[3]\, 
        \MemorySynchronizer_0/SynchStatusReg_168[2]\, 
        \MemorySynchronizer_0/SynchStatusReg_168[1]\, 
        \MemorySynchronizer_0/SynchStatusReg_168[0]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[31]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[30]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[29]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[28]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[27]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[26]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[25]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[24]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[23]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[22]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[21]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[20]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[19]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[18]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[17]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[16]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[15]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[14]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[13]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[12]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[11]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[10]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[9]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[8]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[7]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[6]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[5]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[4]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[3]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[2]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[1]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[0]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[31]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[30]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[29]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[28]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[27]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[26]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[25]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[24]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[23]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[22]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[21]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[20]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[19]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[18]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[17]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[16]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[15]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[14]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[13]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[12]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[11]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[10]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[9]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[8]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[7]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[6]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[5]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[4]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[3]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[2]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[1]\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[0]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[31]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[30]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[29]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[28]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[27]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[26]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[25]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[24]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[23]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[22]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[21]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[20]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[19]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[18]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[17]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[16]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[15]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[14]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[13]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[12]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[11]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[10]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[9]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[8]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[7]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[6]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[5]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[4]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[3]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[2]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[1]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[0]\, 
        \MemorySynchronizer_0/end_one_counter_Z[1]\, 
        \MemorySynchronizer_0/end_one_counter_Z[0]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[31]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[30]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[29]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[28]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[27]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[26]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[25]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[24]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[23]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[22]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[21]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[20]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[19]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[18]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[17]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[16]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[15]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[14]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[13]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[12]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[11]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[10]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[9]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[8]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[7]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[6]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[5]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[4]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[3]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[2]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[1]\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[0]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_Z[31]\, 
        \MemorySynchronizer_0/numberofpendingresyncrequest_Z[2]\, 
        \MemorySynchronizer_0/numberofpendingresyncrequest_Z[1]\, 
        \MemorySynchronizer_0/numberofpendingresyncrequest_Z[0]\, 
        \MemorySynchronizer_0/ConfigReg_Z[31]\, 
        \MemorySynchronizer_0/ConfigReg_Z[30]\, 
        \MemorySynchronizer_0/ConfigReg_Z[29]\, 
        \MemorySynchronizer_0/ConfigReg_Z[28]\, 
        \MemorySynchronizer_0/ConfigReg_Z[27]\, 
        \MemorySynchronizer_0/ConfigReg_Z[26]\, 
        \MemorySynchronizer_0/ConfigReg_Z[25]\, 
        \MemorySynchronizer_0/ConfigReg_Z[24]\, 
        \MemorySynchronizer_0/ConfigReg_Z[23]\, 
        \MemorySynchronizer_0/ConfigReg_Z[22]\, 
        \MemorySynchronizer_0/ConfigReg_Z[21]\, 
        \MemorySynchronizer_0/ConfigReg_Z[20]\, 
        \MemorySynchronizer_0/ConfigReg_Z[19]\, 
        \MemorySynchronizer_0/ConfigReg_Z[18]\, 
        \MemorySynchronizer_0/ConfigReg_Z[17]\, 
        \MemorySynchronizer_0/ConfigReg_Z[16]\, 
        \MemorySynchronizer_0/ConfigReg_Z[15]\, 
        \MemorySynchronizer_0/ConfigReg_Z[14]\, 
        \MemorySynchronizer_0/ConfigReg_Z[13]\, 
        \MemorySynchronizer_0/ConfigReg_Z[12]\, 
        \MemorySynchronizer_0/ConfigReg_Z[11]\, 
        \MemorySynchronizer_0/ConfigReg_Z[10]\, 
        \MemorySynchronizer_0/ConfigReg_Z[9]\, 
        \MemorySynchronizer_0/ConfigReg_Z[8]\, 
        \MemorySynchronizer_0/ConfigReg_Z[7]\, 
        \MemorySynchronizer_0/ConfigReg_Z[6]\, 
        \MemorySynchronizer_0/ConfigReg_Z[5]\, 
        \MemorySynchronizer_0/ConfigReg_Z[4]\, 
        \MemorySynchronizer_0/ConfigReg_Z[3]\, 
        \MemorySynchronizer_0/ConfigReg_Z[2]\, 
        \MemorySynchronizer_0/ConfigReg_Z[1]\, 
        \MemorySynchronizer_0/ConfigReg_Z[0]\, 
        \MemorySynchronizer_0/numberofnewavails_Z[2]\, 
        \MemorySynchronizer_0/numberofnewavails_Z[1]\, 
        \MemorySynchronizer_0/numberofnewavails_Z[0]\, 
        \MemorySynchronizer_0/MemorySyncState_Z[5]\, 
        \MemorySynchronizer_0/MemorySyncState_Z[4]\, 
        \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        \MemorySynchronizer_0/MemorySyncState_Z[2]\, 
        \MemorySynchronizer_0/MemorySyncState_Z[1]\, 
        \MemorySynchronizer_0/MemorySyncState_Z[0]\, 
        \MemorySynchronizer_0/MemorySyncState_ns[4]\, 
        \MemorySynchronizer_0/MemorySyncState_ns[2]\, 
        \MemorySynchronizer_0/MemorySyncState_ns[1]\, 
        \MemorySynchronizer_0/MemorySyncState_ns[0]\, 
        \MemorySynchronizer_0/APBState_ns[1]\, 
        \MemorySynchronizer_0/APBState_ns[0]\, 
        \MemorySynchronizer_0/MemorySyncStatece_Z[0]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[30]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[29]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[28]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[27]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[26]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[25]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[24]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[23]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[22]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[21]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[20]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[19]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[18]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[17]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[16]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[15]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[14]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[13]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[12]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[11]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[10]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[9]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[8]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[7]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[6]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[5]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[4]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[3]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[2]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[1]\, 
        \MemorySynchronizer_0/waitingtimercounterrs[0]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[30]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[29]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[28]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[27]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[26]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[25]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[24]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[23]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[22]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[21]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[20]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[19]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[18]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[17]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[16]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[15]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[14]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[13]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[12]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[11]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[10]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[9]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[8]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[7]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[6]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[5]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[4]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[3]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[2]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[1]\, 
        \MemorySynchronizer_0/waitingtimercounter_Z[0]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[31]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[30]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[29]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[28]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[27]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[26]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[25]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[24]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[23]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[22]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[21]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[20]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[19]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[18]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[17]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[16]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[15]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[14]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[13]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[12]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[11]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[10]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[9]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[8]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[7]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[6]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[5]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[4]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[3]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[2]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[1]\, 
        \MemorySynchronizer_0/waitingtimercounter_10[0]\, 
        \MemorySynchronizer_0/resettimercounterrs[30]\, 
        \MemorySynchronizer_0/resettimercounterrs[29]\, 
        \MemorySynchronizer_0/resettimercounterrs[28]\, 
        \MemorySynchronizer_0/resettimercounterrs[27]\, 
        \MemorySynchronizer_0/resettimercounterrs[26]\, 
        \MemorySynchronizer_0/resettimercounterrs[25]\, 
        \MemorySynchronizer_0/resettimercounterrs[24]\, 
        \MemorySynchronizer_0/resettimercounterrs[23]\, 
        \MemorySynchronizer_0/resettimercounterrs[22]\, 
        \MemorySynchronizer_0/resettimercounterrs[21]\, 
        \MemorySynchronizer_0/resettimercounterrs[20]\, 
        \MemorySynchronizer_0/resettimercounterrs[19]\, 
        \MemorySynchronizer_0/resettimercounterrs[18]\, 
        \MemorySynchronizer_0/resettimercounterrs[17]\, 
        \MemorySynchronizer_0/resettimercounterrs[16]\, 
        \MemorySynchronizer_0/resettimercounterrs[15]\, 
        \MemorySynchronizer_0/resettimercounterrs[14]\, 
        \MemorySynchronizer_0/resettimercounterrs[13]\, 
        \MemorySynchronizer_0/resettimercounterrs[12]\, 
        \MemorySynchronizer_0/resettimercounterrs[11]\, 
        \MemorySynchronizer_0/resettimercounterrs[10]\, 
        \MemorySynchronizer_0/resettimercounterrs[9]\, 
        \MemorySynchronizer_0/resettimercounterrs[8]\, 
        \MemorySynchronizer_0/resettimercounterrs[7]\, 
        \MemorySynchronizer_0/resettimercounterrs[6]\, 
        \MemorySynchronizer_0/resettimercounterrs[5]\, 
        \MemorySynchronizer_0/resettimercounterrs[4]\, 
        \MemorySynchronizer_0/resettimercounterrs[3]\, 
        \MemorySynchronizer_0/resettimercounterrs[2]\, 
        \MemorySynchronizer_0/resettimercounterrs[1]\, 
        \MemorySynchronizer_0/resettimercounterrs[0]\, 
        \MemorySynchronizer_0/resettimercounter_Z[31]\, 
        \MemorySynchronizer_0/resettimercounter_Z[30]\, 
        \MemorySynchronizer_0/resettimercounter_Z[29]\, 
        \MemorySynchronizer_0/resettimercounter_Z[28]\, 
        \MemorySynchronizer_0/resettimercounter_Z[27]\, 
        \MemorySynchronizer_0/resettimercounter_Z[26]\, 
        \MemorySynchronizer_0/resettimercounter_Z[25]\, 
        \MemorySynchronizer_0/resettimercounter_Z[24]\, 
        \MemorySynchronizer_0/resettimercounter_Z[23]\, 
        \MemorySynchronizer_0/resettimercounter_Z[22]\, 
        \MemorySynchronizer_0/resettimercounter_Z[21]\, 
        \MemorySynchronizer_0/resettimercounter_Z[20]\, 
        \MemorySynchronizer_0/resettimercounter_Z[19]\, 
        \MemorySynchronizer_0/resettimercounter_Z[18]\, 
        \MemorySynchronizer_0/resettimercounter_Z[17]\, 
        \MemorySynchronizer_0/resettimercounter_Z[16]\, 
        \MemorySynchronizer_0/resettimercounter_Z[15]\, 
        \MemorySynchronizer_0/resettimercounter_Z[14]\, 
        \MemorySynchronizer_0/resettimercounter_Z[13]\, 
        \MemorySynchronizer_0/resettimercounter_Z[12]\, 
        \MemorySynchronizer_0/resettimercounter_Z[11]\, 
        \MemorySynchronizer_0/resettimercounter_Z[10]\, 
        \MemorySynchronizer_0/resettimercounter_Z[9]\, 
        \MemorySynchronizer_0/resettimercounter_Z[8]\, 
        \MemorySynchronizer_0/resettimercounter_Z[7]\, 
        \MemorySynchronizer_0/resettimercounter_Z[6]\, 
        \MemorySynchronizer_0/resettimercounter_Z[5]\, 
        \MemorySynchronizer_0/resettimercounter_Z[4]\, 
        \MemorySynchronizer_0/resettimercounter_Z[3]\, 
        \MemorySynchronizer_0/resettimercounter_Z[2]\, 
        \MemorySynchronizer_0/resettimercounter_Z[1]\, 
        \MemorySynchronizer_0/resettimercounter_Z[0]\, 
        \MemorySynchronizer_0/resettimercounter_9[31]\, 
        \MemorySynchronizer_0/resettimercounter_9[30]\, 
        \MemorySynchronizer_0/resettimercounter_9[29]\, 
        \MemorySynchronizer_0/resettimercounter_9[28]\, 
        \MemorySynchronizer_0/resettimercounter_9[27]\, 
        \MemorySynchronizer_0/resettimercounter_9[26]\, 
        \MemorySynchronizer_0/resettimercounter_9[25]\, 
        \MemorySynchronizer_0/resettimercounter_9[24]\, 
        \MemorySynchronizer_0/resettimercounter_9[23]\, 
        \MemorySynchronizer_0/resettimercounter_9[22]\, 
        \MemorySynchronizer_0/resettimercounter_9[21]\, 
        \MemorySynchronizer_0/resettimercounter_9[20]\, 
        \MemorySynchronizer_0/resettimercounter_9[19]\, 
        \MemorySynchronizer_0/resettimercounter_9[18]\, 
        \MemorySynchronizer_0/resettimercounter_9[17]\, 
        \MemorySynchronizer_0/resettimercounter_9[16]\, 
        \MemorySynchronizer_0/resettimercounter_9[15]\, 
        \MemorySynchronizer_0/resettimercounter_9[14]\, 
        \MemorySynchronizer_0/resettimercounter_9[13]\, 
        \MemorySynchronizer_0/resettimercounter_9[12]\, 
        \MemorySynchronizer_0/resettimercounter_9[11]\, 
        \MemorySynchronizer_0/resettimercounter_9[10]\, 
        \MemorySynchronizer_0/resettimercounter_9[9]\, 
        \MemorySynchronizer_0/resettimercounter_9[8]\, 
        \MemorySynchronizer_0/resettimercounter_9[7]\, 
        \MemorySynchronizer_0/resettimercounter_9[6]\, 
        \MemorySynchronizer_0/resettimercounter_9[5]\, 
        \MemorySynchronizer_0/resettimercounter_9[4]\, 
        \MemorySynchronizer_0/resettimercounter_9[3]\, 
        \MemorySynchronizer_0/resettimercounter_9[2]\, 
        \MemorySynchronizer_0/resettimercounter_9[1]\, 
        \MemorySynchronizer_0/resettimercounter_9[0]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[22]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[21]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[20]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[19]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[18]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[17]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[16]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[15]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[14]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[13]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[12]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[11]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[10]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[9]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[8]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[7]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[6]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[5]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[4]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[3]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[2]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[1]\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[0]\, 
        \MemorySynchronizer_0/resynctimercounter_1[31]\, 
        \MemorySynchronizer_0/resynctimercounter_1[30]\, 
        \MemorySynchronizer_0/resynctimercounter_1[29]\, 
        \MemorySynchronizer_0/resynctimercounter_1[28]\, 
        \MemorySynchronizer_0/resynctimercounter_1[27]\, 
        \MemorySynchronizer_0/resynctimercounter_1[26]\, 
        \MemorySynchronizer_0/resynctimercounter_1[25]\, 
        \MemorySynchronizer_0/resynctimercounter_1[24]\, 
        \MemorySynchronizer_0/resynctimercounter_1[23]\, 
        \MemorySynchronizer_0/resynctimercounter_1[22]\, 
        \MemorySynchronizer_0/resynctimercounter_1[21]\, 
        \MemorySynchronizer_0/resynctimercounter_1[20]\, 
        \MemorySynchronizer_0/resynctimercounter_1[19]\, 
        \MemorySynchronizer_0/resynctimercounter_1[18]\, 
        \MemorySynchronizer_0/resynctimercounter_1[17]\, 
        \MemorySynchronizer_0/resynctimercounter_1[16]\, 
        \MemorySynchronizer_0/resynctimercounter_1[15]\, 
        \MemorySynchronizer_0/resynctimercounter_1[14]\, 
        \MemorySynchronizer_0/resynctimercounter_1[13]\, 
        \MemorySynchronizer_0/resynctimercounter_1[12]\, 
        \MemorySynchronizer_0/resynctimercounter_1[11]\, 
        \MemorySynchronizer_0/resynctimercounter_1[10]\, 
        \MemorySynchronizer_0/resynctimercounter_1[9]\, 
        \MemorySynchronizer_0/resynctimercounter_1[8]\, 
        \MemorySynchronizer_0/resynctimercounter_1[7]\, 
        \MemorySynchronizer_0/resynctimercounter_1[6]\, 
        \MemorySynchronizer_0/resynctimercounter_1[5]\, 
        \MemorySynchronizer_0/resynctimercounter_1[4]\, 
        \MemorySynchronizer_0/resynctimercounter_1[3]\, 
        \MemorySynchronizer_0/resynctimercounter_1[2]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[14]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[13]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[12]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[11]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[10]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[9]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[8]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[7]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[6]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[5]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[4]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[3]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[2]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[1]\, 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[0]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[30]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[29]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[28]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[27]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[26]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[25]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[24]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[23]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[22]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[21]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[20]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[19]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[18]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[17]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[16]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[15]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[14]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[13]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[12]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[11]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[10]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[9]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[8]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[7]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[6]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[5]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[4]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[3]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[2]\, 
        \MemorySynchronizer_0/un120_in_enable_i_A[1]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[30]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[29]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[28]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[27]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[26]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[25]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[24]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[23]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[22]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[21]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[20]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[19]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[18]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[17]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[16]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[15]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[14]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[13]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[12]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[11]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[10]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[9]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[8]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[7]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[6]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[5]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[4]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[3]\, 
        \MemorySynchronizer_0/un120_in_enable_a_4[2]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[15]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[14]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[13]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[12]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[11]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[10]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[9]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[8]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[7]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[6]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[5]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[4]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[3]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[2]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[1]\, 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[0]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_o2_1_0[4]\, 
        \MemorySynchronizer_0/numberofnewavails_RNIVL541_1_Z[0]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_0_0_0[4]\, 
        \MemorySynchronizer_0/SynchStatusReg_RNO_2_Z[5]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_16_0_Z[28]\, 
        \MemorySynchronizer_0/numberofnewavails_RNIEAMF1_Z[0]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_34_1[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_1_1_Z[4]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_31_Z[20]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[26]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[25]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[24]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[23]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[22]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[21]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[20]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[11]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[3]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[2]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[0]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[30]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[29]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[28]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[27]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[26]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[25]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[24]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[23]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[22]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[21]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[20]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[19]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[18]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[17]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[15]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[14]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[12]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[11]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[4]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[3]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[2]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[1]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[0]\, 
        \MemorySynchronizer_0/MemorySyncState_ns_0_0_0_1_Z[4]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_1_Z[11]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_a2_0_Z[1]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_a2_0_Z[0]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_14_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_10_Z[20]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_m_0_0[13]\, 
        \MemorySynchronizer_0/ResetTimerValueReg_m_0_0[6]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_18_0_Z[19]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_2_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_21_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_19_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_18_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_17_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_16_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_15_Z[20]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_0_Z[28]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_Z[28]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_2_0_Z[4]\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[14]\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[12]\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[4]\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[1]\, 
        \MemorySynchronizer_0/SynchStatusReg_m[7]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[29]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[28]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[26]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[25]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[24]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[23]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[22]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[21]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[20]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[18]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[16]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[14]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[13]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[12]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[11]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[10]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[9]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[8]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[7]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[6]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[5]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[4]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[2]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[1]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[0]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_0_Z[15]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_0_Z[3]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[30]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[27]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[19]\, 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[17]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[30]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[29]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[28]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[27]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[26]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[25]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[24]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[22]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[20]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[19]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[17]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[16]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[14]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[13]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[10]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[9]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[6]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[4]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[2]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[1]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[0]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_25_Z[20]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[32]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[31]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[30]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[28]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[23]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[22]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[18]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[16]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[15]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[13]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[12]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[10]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[8]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[7]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[6]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[5]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[4]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[3]\, 
        \MemorySynchronizer_0/un5_resettimercounter_m[2]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_28_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_27_Z[20]\, 
        \MemorySynchronizer_0/MemorySyncState_ns_0_0_Z[1]\, 
        \MemorySynchronizer_0/MemorySyncState_ns_0_1_Z[0]\, 
        \MemorySynchronizer_0/resettimercounter_m[13]\, 
        \MemorySynchronizer_0/resettimercounter_m[6]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_0_Z[4]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[23]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[21]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[18]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[15]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[12]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[11]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[8]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[7]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[5]\, 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[3]\, 
        \MemorySynchronizer_0/SynchStatusReg_152_Z[30]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[30]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[28]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[16]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[13]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[9]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[8]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[6]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[4]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[1]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[31]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[30]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[29]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[28]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[27]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[26]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[25]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[24]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[23]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[22]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[21]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[20]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[19]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[18]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[17]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[15]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[14]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[12]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[11]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[10]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[9]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[7]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[5]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[4]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[3]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[2]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[1]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[0]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[31]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[29]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[27]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[26]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[25]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[24]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[23]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[22]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[21]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[20]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[19]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[18]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[17]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[16]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[15]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[14]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[13]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[12]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[11]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[10]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[9]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[8]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[7]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[6]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[5]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[3]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[2]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[0]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_1_0[7]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[10]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[31]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[30]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[29]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[28]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[27]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[19]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[18]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[17]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[16]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[15]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[14]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[13]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[12]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[8]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[6]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[5]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[4]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[1]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[16]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[13]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[10]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[9]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[8]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[7]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[6]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[26]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[25]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[24]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[23]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[22]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[21]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[20]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[11]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[3]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[2]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[0]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[31]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[10]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[9]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[7]\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[5]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_0_a2_0_0_Z[25]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_0_a2_0_0_Z[22]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_2_0_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_4_0_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_3_0_Z[20]\, 
        \MemorySynchronizer_0/SynchStatusReg_82_m[5]\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_57_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_58_Z\, 
        \MemorySynchronizer_0/N_1978_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_51_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_52_i_i_a2_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_53_i_i_a2_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_40_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_41_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_42_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_43_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_44_Z\, 
        \MemorySynchronizer_0/N_1979_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_35_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_59_Z\, 
        \MemorySynchronizer_0/N_1981_i\, 
        \MemorySynchronizer_0/N_21_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_60_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_54_i_i_a2_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_33_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_46_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_56_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_36_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_34_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_32_i_i_a2_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_55_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_47_i_i_a2_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_48_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_49_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_37_Z\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_38_Z\, 
        \MemorySynchronizer_0/N_1980_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_52\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_53\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_54\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_55\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_56_i_i_a2_Z\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_57_i_i_a2_Z\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_58_i_i_a2_Z\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_59\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_60\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_36\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_41\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_48\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_34\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_49\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_47\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_43\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_44\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_45\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_46\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_51\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_50\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_37\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_40\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_39\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_32\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_31\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_35\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_61\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_33\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_38\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_42\, 
        \MemorySynchronizer_0/temp_1_cry_0_Y\, 
        \MemorySynchronizer_0/N_1158_i_i\, 
        \MemorySynchronizer_0/N_527_i_i\, 
        \MemorySynchronizer_0/N_1052_i_i\, 
        \MemorySynchronizer_0/N_2032_i\, 
        \MemorySynchronizer_0/N_215_i\, 
        \MemorySynchronizer_0/N_2033_i\, 
        \MemorySynchronizer_0/N_2034_i\, 
        \MemorySynchronizer_0/N_2035_i\, 
        \MemorySynchronizer_0/SynchStatusReg_152_e2\, 
        \MemorySynchronizer_0/N_113_i\, 
        \MemorySynchronizer_0/N_2015_i\, 
        \MemorySynchronizer_0/N_2016_i\, 
        \MemorySynchronizer_0/N_1104\, 
        \MemorySynchronizer_0/N_699\, 
        \MemorySynchronizer_0/N_1103\, 
        \MemorySynchronizer_0/N_1102\, 
        \MemorySynchronizer_0/N_1101\, 
        \MemorySynchronizer_0/N_1100\, 
        \MemorySynchronizer_0/N_1099\, 
        \MemorySynchronizer_0/N_1098\, 
        \MemorySynchronizer_0/N_1097\, 
        \MemorySynchronizer_0/N_1096\, 
        \MemorySynchronizer_0/N_1095\, 
        \MemorySynchronizer_0/N_1094\, 
        \MemorySynchronizer_0/N_1093\, 
        \MemorySynchronizer_0/N_1092\, 
        \MemorySynchronizer_0/N_1119\, 
        \MemorySynchronizer_0/N_1118\, 
        \MemorySynchronizer_0/N_1117\, 
        \MemorySynchronizer_0/N_1116\, 
        \MemorySynchronizer_0/N_1115\, 
        \MemorySynchronizer_0/N_1114\, 
        \MemorySynchronizer_0/N_1113\, 
        \MemorySynchronizer_0/N_1112\, 
        \MemorySynchronizer_0/N_1111\, 
        \MemorySynchronizer_0/N_1110\, 
        \MemorySynchronizer_0/N_1109\, 
        \MemorySynchronizer_0/N_1108\, 
        \MemorySynchronizer_0/N_1107\, 
        \MemorySynchronizer_0/N_1106\, 
        \MemorySynchronizer_0/N_1105\, 
        \MemorySynchronizer_0/N_1122\, 
        \MemorySynchronizer_0/N_1121\, 
        \MemorySynchronizer_0/N_1120\, 
        \MemorySynchronizer_0/N_2304_i\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_Z\, 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0_Z\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, 
        \MemorySynchronizer_0/N_207_i\, 
        \MemorySynchronizer_0/N_2030_i\, 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, 
        \MemorySynchronizer_0/un104_in_enable_16\, 
        \MemorySynchronizer_0/un104_in_enable_17\, 
        \MemorySynchronizer_0/un104_in_enable_18\, 
        \MemorySynchronizer_0/un104_in_enable_19\, 
        \MemorySynchronizer_0/un104_in_enable_20\, 
        \MemorySynchronizer_0/un104_in_enable_21\, 
        \MemorySynchronizer_0/un104_in_enable_22\, 
        \MemorySynchronizer_0/un104_in_enable_23\, 
        \MemorySynchronizer_0/un104_in_enable_24\, 
        \MemorySynchronizer_0/un104_in_enable_25\, 
        \MemorySynchronizer_0/un104_in_enable_26\, 
        \MemorySynchronizer_0/un104_in_enable_27\, 
        \MemorySynchronizer_0/un104_in_enable_28\, 
        \MemorySynchronizer_0/un104_in_enable_29\, 
        \MemorySynchronizer_0/un104_in_enable_30\, 
        \MemorySynchronizer_0/un104_in_enable_1\, 
        \MemorySynchronizer_0/un104_in_enable_2\, 
        \MemorySynchronizer_0/un104_in_enable_3\, 
        \MemorySynchronizer_0/un104_in_enable_4\, 
        \MemorySynchronizer_0/un104_in_enable_5\, 
        \MemorySynchronizer_0/un104_in_enable_6\, 
        \MemorySynchronizer_0/un104_in_enable_7\, 
        \MemorySynchronizer_0/un104_in_enable_8\, 
        \MemorySynchronizer_0/un104_in_enable_9\, 
        \MemorySynchronizer_0/un104_in_enable_10\, 
        \MemorySynchronizer_0/un104_in_enable_11\, 
        \MemorySynchronizer_0/un104_in_enable_12\, 
        \MemorySynchronizer_0/un104_in_enable_13\, 
        \MemorySynchronizer_0/un104_in_enable_14\, 
        \MemorySynchronizer_0/un104_in_enable_15\, 
        \MemorySynchronizer_0/un104_in_enable_0\, 
        \MemorySynchronizer_0/numberofnewavails_0_sqmuxa\, 
        \MemorySynchronizer_0/ConfigReg_0\, 
        \MemorySynchronizer_0/N_2305_i\, 
        \MemorySynchronizer_0/un1_APBState_i\, 
        \MemorySynchronizer_0/N_2306_i\, 
        \MemorySynchronizer_0/N_304\, 
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa_i\, 
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa_1_i_Z\, 
        \MemorySynchronizer_0/N_191_i\, 
        \MemorySynchronizer_0/ReadInterrupt_0_sqmuxa_2_i_0_0_Z\, 
        \MemorySynchronizer_0/N_2068_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_42_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_35_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_35_i\, 
        \MemorySynchronizer_0/un104_in_enable_axb_31\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_38_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_51_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_51_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_33_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_47_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_47_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_61_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_24_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_24_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_35_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_46_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_46_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_31_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_40_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_40_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_32_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_62_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_62_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_39_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_43_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_43_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_40_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_22_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_22_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_37_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_25_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_25_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_50_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_42_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_42_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_51_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_26_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_26_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_46_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_39_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_39_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_45_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_38_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_38_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_44_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_37_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_37_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_43_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_36_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_36_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_47_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_20_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_20_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_49_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_1_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_1_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_34_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_45_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_45_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_48_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_2_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_2_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_41_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_4_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_4_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_36_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_5_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_5_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_60_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_60_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_60_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_59_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_59_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_59_i\, 
        \MemorySynchronizer_0/N_2532_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_58_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_58_i\, 
        \MemorySynchronizer_0/N_2533_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_57_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_57_i\, 
        \MemorySynchronizer_0/N_2534_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_56_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_56_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_55_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_55_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_55_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_54_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_54_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_54_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_53_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_53_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_53_i\, 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_52_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_52_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_52_i\, 
        \MemorySynchronizer_0/N_1980_i_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_12_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_12_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_38_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_11_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_11_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_37_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_10_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_10_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_49_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_9_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_9_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_48_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_29_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_29_i\, 
        \MemorySynchronizer_0/N_2538_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_28_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_28_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_55_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_27_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_27_i\, 
        \MemorySynchronizer_0/N_2539_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_19_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_19_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_34_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_8_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_8_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_36_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_6_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_6_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_56_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_49_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_49_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_46_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_48_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_48_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_33_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_61_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_61_i\, 
        \MemorySynchronizer_0/N_2535_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_44_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_44_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_60_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_23_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_23_i\, 
        \MemorySynchronizer_0/N_21_i_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_3_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_3_i\, 
        \MemorySynchronizer_0/N_1981_i_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_41_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_41_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_59_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_21_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_21_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_35_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_7_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_7_i\, 
        \MemorySynchronizer_0/N_1979_i_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_18_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_18_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_44_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_17_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_17_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_43_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_16_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_16_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_42_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_15_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_15_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_41_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_14_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_14_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_40_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_13_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_13_i\, 
        \MemorySynchronizer_0/N_2536_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_34_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_34_i\, 
        \MemorySynchronizer_0/N_2537_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_33_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_33_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_51_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_32_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_32_i\, 
        \MemorySynchronizer_0/N_1978_i_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_31_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_31_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_58_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_30_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_30_i\, 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_57_set_Z\, 
        \MemorySynchronizer_0/un1_nreset_50_rs_Z\, 
        \MemorySynchronizer_0/un1_nreset_50_i\, 
        \MemorySynchronizer_0/N_301\, 
        \MemorySynchronizer_0/enableTimestampGen_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_0_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_1_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_1_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_2_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_2_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_3_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_3_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_4_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_4_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_5_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_5_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_6_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_6_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_7_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_7_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_8_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_8_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_9_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_9_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_10_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_10_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_11_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_11_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_12_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_12_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_13_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_13_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_14_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_14_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_15_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_15_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_16_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_16_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_17_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_17_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_18_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_18_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_19_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_19_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_20_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_20_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_21_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_21_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_22_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_22_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_23_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_23_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_24_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_24_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_25_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_25_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_26_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_26_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_27_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_27_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_28_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_28_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_29_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_29_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_s_31_S\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_30_Z\, 
        \MemorySynchronizer_0/un5_resettimercounter_cry_30_S\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_0_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_1_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_2_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_3_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_4_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_5_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_6_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_7_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_8_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_9_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_10_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_11_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_12_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_13_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_14_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_15_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_16_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_17_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_18_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_19_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_20_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_21_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_22_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_23_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_24_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_25_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_26_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_27_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_28_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_29_Z\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, 
        \MemorySynchronizer_0/temp_1_cry_0\, 
        \MemorySynchronizer_0/temp_1_cry_1\, 
        \MemorySynchronizer_0/temp_1_cry_2\, 
        \MemorySynchronizer_0/temp_1_cry_3\, 
        \MemorySynchronizer_0/temp_1_cry_4\, 
        \MemorySynchronizer_0/temp_1_cry_5\, 
        \MemorySynchronizer_0/temp_1_cry_6\, 
        \MemorySynchronizer_0/temp_1_cry_7\, 
        \MemorySynchronizer_0/temp_1_cry_8\, 
        \MemorySynchronizer_0/temp_1_cry_9\, 
        \MemorySynchronizer_0/temp_1_cry_10\, 
        \MemorySynchronizer_0/temp_1_cry_11\, 
        \MemorySynchronizer_0/temp_1_cry_12\, 
        \MemorySynchronizer_0/temp_1_cry_13\, 
        \MemorySynchronizer_0/temp_1_cry_14\, 
        \MemorySynchronizer_0/temp_1_cry_15\, 
        \MemorySynchronizer_0/temp_1_cry_16\, 
        \MemorySynchronizer_0/temp_1_cry_17\, 
        \MemorySynchronizer_0/temp_1_cry_18\, 
        \MemorySynchronizer_0/temp_1_cry_19\, 
        \MemorySynchronizer_0/temp_1_cry_20\, 
        \MemorySynchronizer_0/temp_1_cry_21\, 
        \MemorySynchronizer_0/temp_1_cry_22\, 
        \MemorySynchronizer_0/temp_1_cry_23\, 
        \MemorySynchronizer_0/temp_1_cry_24\, 
        \MemorySynchronizer_0/temp_1_cry_25\, 
        \MemorySynchronizer_0/temp_1_cry_26\, 
        \MemorySynchronizer_0/temp_1_cry_27\, 
        \MemorySynchronizer_0/temp_1_cry_28\, 
        \MemorySynchronizer_0/temp_1_cry_29\, 
        \MemorySynchronizer_0/temp_1_cry_30\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0_Y\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_Y\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_1_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_1_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_2_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_2_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_3_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_3_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_4_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_4_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_5_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_5_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_6_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_6_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_7_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_7_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_8_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_8_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_9_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_9_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_10_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_10_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_11_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_11_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_12_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_12_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_13_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_13_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_14_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_14_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_15_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_15_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_16_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_16_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_17_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_17_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_18_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_18_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_19_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_19_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_20_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_20_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_21_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_21_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_22_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_22_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_23_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_23_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_24_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_24_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_25_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_25_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_26_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_26_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_27_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_27_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_28_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_28_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_29_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_29_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_s_31_S\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_30_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_30_S\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, 
        \MemorySynchronizer_0/un105_m1_e_0_0\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_1_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_2_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_3_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_4_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_5_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_6_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_7_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_8_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_9_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_10_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_11_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_12_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_13_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_14_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_15_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_16_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_17_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_18_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_19_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_20_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_21_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_22_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_23_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_24_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_25_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_26_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_27_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_28_Z\, 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_29_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_0_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_1_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_2_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_3_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_4_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_5_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_6_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_7_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_8_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_9_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_10_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_11_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_12_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_13_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_14_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_15_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_16_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_17_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_18_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_19_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_20_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_21_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_22_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_23_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_24_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_25_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_26_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_27_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_28_Z\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_0_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_1_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_2_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_3_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_4_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_5_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_6_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_7_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_8_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_9_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_10_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_11_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_12_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_13_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_14_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_15_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_16_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_17_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_18_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_19_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_20_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_21_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_22_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_23_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_24_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_25_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_26_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_27_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_28_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_29_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_30_Z\, 
        \MemorySynchronizer_0/un104_in_enable_cry_31_Z\, 
        \MemorySynchronizer_0/un1_in_enable_2_0_0_a2_0_Z\, 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1_0_a2_1_Z\, 
        \MemorySynchronizer_0/N_1076\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_7_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_21_x_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_20_x_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2_N_2L1_1_Z\, 
        \MemorySynchronizer_0/N_2313\, 
        \MemorySynchronizer_0/N_140_1_i\, 
        \MemorySynchronizer_0/N_140_2\, 
        \MemorySynchronizer_0/N_2326\, 
        \MemorySynchronizer_0/N_140_i_1\, 
        \MemorySynchronizer_0/N_140_i\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_28_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_29_Z\, 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa_i_1_i_a2_1_Z\, 
        \MemorySynchronizer_0/N_271\, 
        \MemorySynchronizer_0/N_2569\, \MemorySynchronizer_0/N_6\, 
        \MemorySynchronizer_0/un112_in_enable_0_I_45_RNIRI17A_Z\, 
        \MemorySynchronizer_0/g1\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_22_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_23_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2_1\, 
        \MemorySynchronizer_0/N_2330\, \MemorySynchronizer_0/N_4\, 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_N_2L1_Z\, 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa_i_0_i_a2_1_Z\, 
        \MemorySynchronizer_0/g2_0_0\, 
        \MemorySynchronizer_0/N_2606\, 
        \MemorySynchronizer_0/m3_e_0_0\, 
        \MemorySynchronizer_0/g3\, 
        \MemorySynchronizer_0/N_2028_i\, 
        \MemorySynchronizer_0/SynchStatusReg_2_sqmuxa_1\, 
        \MemorySynchronizer_0/g0_0_1\, 
        \MemorySynchronizer_0/N_2321\, 
        \MemorySynchronizer_0/N_1512\, 
        \MemorySynchronizer_0/N_2310\, 
        \MemorySynchronizer_0/N_2510\, \MemorySynchronizer_0/g2\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_0_Z\, 
        \MemorySynchronizer_0/SynchStatusReg_N_3_mux\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_1_Z\, 
        \MemorySynchronizer_0/N_2604\, 
        \MemorySynchronizer_0/un1_enabletimestampgen2_2_sn\, 
        \MemorySynchronizer_0/N_2575\, 
        \MemorySynchronizer_0/N_1179\, 
        \MemorySynchronizer_0/N_2585\, 
        \MemorySynchronizer_0/N_2582\, 
        \MemorySynchronizer_0/un151_in_enablelto30_19\, 
        \MemorySynchronizer_0/un151_in_enablelto30_23\, 
        \MemorySynchronizer_0/un151_in_enablelto31_1\, 
        \MemorySynchronizer_0/un151_in_enable\, 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_13_Z\, 
        \MemorySynchronizer_0/N_2564\, 
        \MemorySynchronizer_0/N_2567\, 
        \MemorySynchronizer_0/N_2328\, 
        \MemorySynchronizer_0/N_2333\, 
        \MemorySynchronizer_0/un6_in_enable_i_0\, 
        \MemorySynchronizer_0/N_1495\, 
        \MemorySynchronizer_0/N_1482\, 
        \MemorySynchronizer_0/N_1091\, 
        \MemorySynchronizer_0/N_1061\, 
        \MemorySynchronizer_0/N_1062\, 
        \MemorySynchronizer_0/N_1063\, 
        \MemorySynchronizer_0/N_1064\, 
        \MemorySynchronizer_0/N_1065\, 
        \MemorySynchronizer_0/N_1066\, 
        \MemorySynchronizer_0/N_1067\, 
        \MemorySynchronizer_0/N_1068\, 
        \MemorySynchronizer_0/N_1069\, 
        \MemorySynchronizer_0/N_1070\, 
        \MemorySynchronizer_0/N_1071\, 
        \MemorySynchronizer_0/N_1072\, 
        \MemorySynchronizer_0/N_1073\, 
        \MemorySynchronizer_0/N_1074\, 
        \MemorySynchronizer_0/N_1075\, 
        \MemorySynchronizer_0/N_1077\, 
        \MemorySynchronizer_0/N_1078\, 
        \MemorySynchronizer_0/N_1079\, 
        \MemorySynchronizer_0/N_1080\, 
        \MemorySynchronizer_0/N_1081\, 
        \MemorySynchronizer_0/N_1082\, 
        \MemorySynchronizer_0/N_1083\, 
        \MemorySynchronizer_0/N_1084\, 
        \MemorySynchronizer_0/N_1085\, 
        \MemorySynchronizer_0/N_1086\, 
        \MemorySynchronizer_0/N_1087\, 
        \MemorySynchronizer_0/N_1088\, 
        \MemorySynchronizer_0/N_1089\, 
        \MemorySynchronizer_0/N_1090\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_21_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_20_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_19_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_18_Z\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_17_Z\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_0_a1_1_Z\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a1_0_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a1_0_0_Z\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_1_Z\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_23_Z\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_21_Z\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_20_Z\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_19_Z\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_18_Z\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_17_Z\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_16_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_22_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_21_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_20_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_19_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_17_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_16_Z\, 
        \MemorySynchronizer_0/un151_in_enablelto30_17\, 
        \MemorySynchronizer_0/un151_in_enablelto30_16\, 
        \MemorySynchronizer_0/un151_in_enablelto30_15\, 
        \MemorySynchronizer_0/un151_in_enablelto30_14\, 
        \MemorySynchronizer_0/un151_in_enablelto30_13\, 
        \MemorySynchronizer_0/un94_in_enable_23_Z\, 
        \MemorySynchronizer_0/un94_in_enable_22_Z\, 
        \MemorySynchronizer_0/un94_in_enable_21_Z\, 
        \MemorySynchronizer_0/un94_in_enable_20_Z\, 
        \MemorySynchronizer_0/un94_in_enable_19_Z\, 
        \MemorySynchronizer_0/un94_in_enable_18_Z\, 
        \MemorySynchronizer_0/un94_in_enable_17_Z\, 
        \MemorySynchronizer_0/un94_in_enable_16_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_22_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_21_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_20_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_19_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_18_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_17_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_16_Z\, 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_15_Z\, 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, 
        \MemorySynchronizer_0/N_2439\, 
        \MemorySynchronizer_0/N_2553\, 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, 
        \MemorySynchronizer_0/resettimercounter_0_sqmuxa_1\, 
        \MemorySynchronizer_0/N_1209\, 
        \MemorySynchronizer_0/N_1213\, 
        \MemorySynchronizer_0/N_1474\, 
        \MemorySynchronizer_0/N_1480\, 
        \MemorySynchronizer_0/N_2418\, 
        \MemorySynchronizer_0/N_2422\, 
        \MemorySynchronizer_0/N_1493\, 
        \MemorySynchronizer_0/N_1497\, 
        \MemorySynchronizer_0/N_1501\, 
        \MemorySynchronizer_0/N_1505\, 
        \MemorySynchronizer_0/N_1509\, 
        \MemorySynchronizer_0/N_1513\, 
        \MemorySynchronizer_0/N_1517\, 
        \MemorySynchronizer_0/N_1521\, 
        \MemorySynchronizer_0/N_1525\, 
        \MemorySynchronizer_0/N_1529\, 
        \MemorySynchronizer_0/N_1533\, 
        \MemorySynchronizer_0/N_1537\, 
        \MemorySynchronizer_0/N_1541\, 
        \MemorySynchronizer_0/N_1549\, 
        \MemorySynchronizer_0/N_1553\, 
        \MemorySynchronizer_0/N_1557\, 
        \MemorySynchronizer_0/N_1561\, 
        \MemorySynchronizer_0/N_1565\, 
        \MemorySynchronizer_0/N_2430\, 
        \MemorySynchronizer_0/N_2315\, 
        \MemorySynchronizer_0/N_2471\, 
        \MemorySynchronizer_0/N_1545\, 
        \MemorySynchronizer_0/N_2337\, 
        \MemorySynchronizer_0/N_2434\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_27_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_25_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_23_Z\, 
        \MemorySynchronizer_0/N_2316\, 
        \MemorySynchronizer_0/SynchStatusReg_152_sm0\, 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, 
        \MemorySynchronizer_0/N_88\, \MemorySynchronizer_0/N_84\, 
        \MemorySynchronizer_0/N_80\, \MemorySynchronizer_0/N_76\, 
        \MemorySynchronizer_0/N_72\, \MemorySynchronizer_0/N_68\, 
        \MemorySynchronizer_0/N_64\, \MemorySynchronizer_0/N_60\, 
        \MemorySynchronizer_0/N_56\, \MemorySynchronizer_0/N_52\, 
        \MemorySynchronizer_0/SynchStatusReg_152_ss0_i_0\, 
        \MemorySynchronizer_0/N_122_i\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_25_Z\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_24_Z\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_23_Z\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_22_Z\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_21_Z\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_19_Z\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_18_Z\, 
        \MemorySynchronizer_0/un6_in_enable_0_a3_28_Z\, 
        \MemorySynchronizer_0/un94_in_enable_29_Z\, 
        \MemorySynchronizer_0/un94_in_enable_28_Z\, 
        \MemorySynchronizer_0/N_2317\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_27_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_30_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_29_Z\, 
        \MemorySynchronizer_0/N_2509\, 
        \MemorySynchronizer_0/N_2576\, 
        \MemorySynchronizer_0/N_2595\, 
        \MemorySynchronizer_0/N_2596\, 
        \MemorySynchronizer_0/un41_in_enable_i_0\, 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_0_a1_Z\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a1_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_0_a1_Z\, 
        \MemorySynchronizer_0/N_2561\, 
        \MemorySynchronizer_0/N_2572\, 
        \MemorySynchronizer_0/N_1182\, 
        \MemorySynchronizer_0/N_2580\, 
        \MemorySynchronizer_0/N_2581\, 
        \MemorySynchronizer_0/N_2586\, 
        \MemorySynchronizer_0/N_2598\, 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_31_Z\, 
        \MemorySynchronizer_0/N_2593\, 
        \MemorySynchronizer_0/N_1201\, 
        \MemorySynchronizer_0/N_1365\, 
        \MemorySynchronizer_0/N_2588\, 
        \MemorySynchronizer_0/N_2323\, 
        \MemorySynchronizer_0/N_2597\, 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a0_1_Z\, 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_4_Z\, 
        \MemorySynchronizer_0/N_1163\, 
        \MemorySynchronizer_0/N_1172\, 
        \MemorySynchronizer_0/N_1217\, 
        \MemorySynchronizer_0/N_1228\, 
        \MemorySynchronizer_0/N_1236\, 
        \MemorySynchronizer_0/N_1245\, 
        \MemorySynchronizer_0/N_1254\, 
        \MemorySynchronizer_0/N_2517\, 
        \MemorySynchronizer_0/N_2574\, 
        \MemorySynchronizer_0/N_2577\, 
        \MemorySynchronizer_0/N_2594\, 
        \MemorySynchronizer_0/N_1123\, 
        \MemorySynchronizer_0/N_1204_1\, 
        \MemorySynchronizer_0/N_1260\, 
        \MemorySynchronizer_0/N_1168\, 
        \MemorySynchronizer_0/N_1177\, 
        \MemorySynchronizer_0/N_1222\, 
        \MemorySynchronizer_0/N_1342\, 
        \MemorySynchronizer_0/N_1403\, 
        \MemorySynchronizer_0/N_1411\, 
        \MemorySynchronizer_0/N_1437\, 
        \MemorySynchronizer_0/N_1445\, 
        \MemorySynchronizer_0/N_1453\, 
        \MemorySynchronizer_0/N_1461\, 
        \MemorySynchronizer_0/N_1469\, 
        \MemorySynchronizer_0/N_191\, 
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa\, 
        \MemorySynchronizer_0/N_1265\, 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_16_Z\, 
        \MemorySynchronizer_0/SynchStatusReg_N_7\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[30]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[29]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[28]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[27]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[26]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[25]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[24]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[23]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[22]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[21]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[20]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[19]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[18]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[17]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[16]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[15]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[14]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[13]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[12]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[11]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[10]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[9]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[8]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[7]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[6]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[5]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[4]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[3]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[2]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[1]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s[0]\, 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[5]\, 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[4]\, 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[3]\, 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[2]\, 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[1]\, 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[0]\, 
        \MemorySynchronizer_0/TimeStampGen/prescaler_5_Z[4]\, 
        \MemorySynchronizer_0/TimeStampGen/prescaler_5_Z[3]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s_Z[31]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[30]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[29]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[28]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[27]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[26]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[25]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[24]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[23]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[22]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[21]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[20]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[19]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[18]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[17]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[16]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[15]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[14]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[13]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[12]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[11]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[10]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[9]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[8]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[7]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[6]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[5]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[4]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[3]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[2]\, 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[1]\, 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc5_Z\, 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc0_Z\, 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc1_Z\, 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc2_Z\, 
        \MemorySynchronizer_0/TimeStampGen/countere\, 
        \MemorySynchronizer_0/TimeStampGen/counter_s_387_FCO\, 
        \MemorySynchronizer_0/TimeStampGen/un6_enable_3_Z\, 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_c2\, 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_c4\, 
        ff_to_start_net, \stamp0_spi_temp_cs_obuf/U0/DOUT1\, 
        \stamp0_spi_temp_cs_obuf/U0/DOUT\, 
        \stamp0_spi_temp_cs_obuf/U0/EOUT1\, 
        \stamp0_spi_temp_cs_obuf/U0/EOUT\, 
        \adc_start_obuf/U0/DOUT1\, \adc_start_obuf/U0/DOUT\, 
        \adc_start_obuf/U0/EOUT1\, \adc_start_obuf/U0/EOUT\, 
        \MISO_ibuf/U0/YIN1\, \MISO_ibuf/U0/YIN\, 
        \stamp0_spi_clock_obuf/U0/DOUT1\, 
        \stamp0_spi_clock_obuf/U0/DOUT\, 
        \stamp0_spi_clock_obuf/U0/EOUT1\, 
        \stamp0_spi_clock_obuf/U0/EOUT\, 
        \LED_RECORDING_obuf/U0/DOUT1\, 
        \LED_RECORDING_obuf/U0/DOUT\, 
        \LED_RECORDING_obuf/U0/EOUT1\, 
        \LED_RECORDING_obuf/U0/EOUT\, \SCLK_obuf/U0/DOUT1\, 
        \SCLK_obuf/U0/DOUT\, \SCLK_obuf/U0/EOUT1\, 
        \SCLK_obuf/U0/EOUT\, \nCS1_obuf/U0/DOUT1\, 
        \nCS1_obuf/U0/DOUT\, \nCS1_obuf/U0/EOUT1\, 
        \nCS1_obuf/U0/EOUT\, \nCS2_obuf/U0/DOUT1\, 
        \nCS2_obuf/U0/DOUT\, \nCS2_obuf/U0/EOUT1\, 
        \nCS2_obuf/U0/EOUT\, \adc_clk_obuf/U0/DOUT1\, 
        \adc_clk_obuf/U0/DOUT\, \adc_clk_obuf/U0/EOUT1\, 
        \adc_clk_obuf/U0/EOUT\, \ENABLE_MEMORY_LED_obuf/U0/DOUT1\, 
        \ENABLE_MEMORY_LED_obuf/U0/DOUT\, 
        \ENABLE_MEMORY_LED_obuf/U0/EOUT1\, 
        \ENABLE_MEMORY_LED_obuf/U0/EOUT\, 
        \RXSM_SODS_ibuf/U0/YIN1\, \RXSM_SODS_ibuf/U0/YIN\, 
        \sb_sb_0/CCC_0/CCC_INST/CLK0_net\, 
        \sb_sb_0/CCC_0/CCC_INST/CLK1_net\, 
        \sb_sb_0/CCC_0/CCC_INST/CLK2_net\, 
        \sb_sb_0/CCC_0/CCC_INST/CLK3_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX0_SEL_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX1_SEL_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX2_SEL_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX3_SEL_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX0_HOLD_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX1_HOLD_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX2_HOLD_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX3_HOLD_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX0_ARST_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX1_ARST_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX2_ARST_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX3_ARST_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/PLL_BYPASS_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/PLL_ARST_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/PLL_POWERDOWN_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/GPD0_ARST_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/GPD1_ARST_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/GPD2_ARST_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/GPD3_ARST_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/PRESET_N_net\, 
        \sb_sb_0/CCC_0/CCC_INST/PCLK_net\, 
        \sb_sb_0/CCC_0/CCC_INST/PSEL_net\, 
        \sb_sb_0/CCC_0/CCC_INST/PENABLE_net\, 
        \sb_sb_0/CCC_0/CCC_INST/PWRITE_net\, 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[7]\, 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[6]\, 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[5]\, 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[4]\, 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[3]\, 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[2]\, 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[7]\, 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[6]\, 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[5]\, 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[4]\, 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[3]\, 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[2]\, 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[1]\, 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[0]\, 
        \stamp0_ready_dms1_ibuf/U0/YIN1\, 
        \stamp0_ready_dms1_ibuf/U0/YIN\, 
        \debug_led_obuf/U0/DOUT1\, \debug_led_obuf/U0/DOUT\, 
        \debug_led_obuf/U0/EOUT1\, \debug_led_obuf/U0/EOUT\, 
        \RXSM_SOE_ibuf/U0/YIN1\, \RXSM_SOE_ibuf/U0/YIN\, 
        \stamp0_spi_mosi_obuft/U0/DOUT1\, 
        \stamp0_spi_mosi_obuft/U0/DOUT\, 
        \stamp0_spi_mosi_obuft/U0/EOUT1\, 
        \stamp0_spi_mosi_obuft/U0/EOUT\, 
        \stamp0_spi_dms2_cs_obuf/U0/DOUT1\, 
        \stamp0_spi_dms2_cs_obuf/U0/DOUT\, 
        \stamp0_spi_dms2_cs_obuf/U0/EOUT1\, 
        \stamp0_spi_dms2_cs_obuf/U0/EOUT\, 
        \sb_sb_0/SYSRESET_POR/UTDO_net\, 
        \stamp0_ready_temp_ibuf/U0/YIN1\, 
        \stamp0_ready_temp_ibuf/U0/YIN\, 
        \stamp0_spi_miso_ibuf/U0/YIN1\, 
        \stamp0_spi_miso_ibuf/U0/YIN\, 
        \MMUART_0_TXD_M2F_obuf/U0/DOUT1\, 
        \MMUART_0_TXD_M2F_obuf/U0/DOUT\, 
        \MMUART_0_TXD_M2F_obuf/U0/EOUT1\, 
        \MMUART_0_TXD_M2F_obuf/U0/EOUT\, 
        \LED_HEARTBEAT_obuf/U0/DOUT1\, 
        \LED_HEARTBEAT_obuf/U0/DOUT\, 
        \LED_HEARTBEAT_obuf/U0/EOUT1\, 
        \LED_HEARTBEAT_obuf/U0/EOUT\, \MOSI_obuf/U0/DOUT1\, 
        \MOSI_obuf/U0/DOUT\, \MOSI_obuf/U0/EOUT1\, 
        \MOSI_obuf/U0/EOUT\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/COLF_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CRSF_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2HCALIB_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDIF_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_DVF_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_ERRF_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_EV_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CLK_BASE_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_BREADY_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_RREADY_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WLAST_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WVALID_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0]\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net\, 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PRESET_N_net\, 
        \stamp0_spi_dms1_cs_obuf/U0/DOUT1\, 
        \stamp0_spi_dms1_cs_obuf/U0/DOUT\, 
        \stamp0_spi_dms1_cs_obuf/U0/EOUT1\, 
        \stamp0_spi_dms1_cs_obuf/U0/EOUT\, \resetn_obuf/U0/DOUT1\, 
        \resetn_obuf/U0/DOUT\, \resetn_obuf/U0/EOUT1\, 
        \resetn_obuf/U0/EOUT\, \stamp0_ready_dms2_ibuf/U0/YIN1\, 
        \stamp0_ready_dms2_ibuf/U0/YIN\, \RXSM_LO_ibuf/U0/YIN1\, 
        \RXSM_LO_ibuf/U0/YIN\, \MMUART_0_RXD_F2M_ibuf/U0/YIN1\, 
        \MMUART_0_RXD_F2M_ibuf/U0/YIN\, 
        \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_30_FCNET1\, 
        \MemorySynchronizer_0/un112_in_enable_0_I_45_FCNET1\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_FCNET1\, 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_RNIKHI89_FCNET1\, 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_FCNET1\, 
        \STAMP_0/un45_async_state_cry_5_FCNET1\, 
        \MemorySynchronizer_0/un104_in_enable_cry_31_FCNET1\, 
        CFG0_GND_INST_NET, \AND2_0_RNIKOS1/U0_RGB1_YR\, 
        \AND2_0_RNIKOS1/U0_RGB1_RGB0_rgbr_net_1\, 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, 
        \AND2_0_RNIKOS1/U0_RGB1_RGB5_rgbr_net_1\, 
        \AND2_0_RNIKOS1/U0_RGB1_RGB6_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_YR\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB0_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB1_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_YR\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbl_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB12_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB14_rgbr_net_1\, 
        \sb_sb_0/CCC_0/GL1_INST/U0_RGB1_YR\, 
        \sb_sb_0/CCC_0/GL1_INST/U0_YNn_GSouth\, 
        \ResetAND_RNIMHJB/U0_YNn_GSouth\, 
        \AND2_0_RNIKOS1/U0_YNn_GSouth\, 
        \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ADLIB_GND0, 
        ADLIB_VCC1, CI_TO_CO2, CI_TO_CO3, NET_CC_CONFIG4, 
        NET_CC_CONFIG5, NET_CC_CONFIG6, NET_CC_CONFIG7, 
        NET_CC_CONFIG8, NET_CC_CONFIG9, NET_CC_CONFIG10, 
        NET_CC_CONFIG11, NET_CC_CONFIG12, NET_CC_CONFIG13, 
        NET_CC_CONFIG14, NET_CC_CONFIG15, NET_CC_CONFIG16, 
        NET_CC_CONFIG17, NET_CC_CONFIG18, NET_CC_CONFIG19, 
        NET_CC_CONFIG20, NET_CC_CONFIG21, NET_CC_CONFIG22, 
        NET_CC_CONFIG23, NET_CC_CONFIG24, NET_CC_CONFIG25, 
        NET_CC_CONFIG26, NET_CC_CONFIG27, NET_CC_CONFIG28, 
        NET_CC_CONFIG29, NET_CC_CONFIG30, NET_CC_CONFIG31, 
        NET_CC_CONFIG32, NET_CC_CONFIG33, NET_CC_CONFIG34, 
        NET_CC_CONFIG35, NET_CC_CONFIG36, NET_CC_CONFIG37, 
        NET_CC_CONFIG38, NET_CC_CONFIG39, NET_CC_CONFIG40, 
        NET_CC_CONFIG41, NET_CC_CONFIG42, NET_CC_CONFIG43, 
        NET_CC_CONFIG44, NET_CC_CONFIG45, NET_CC_CONFIG46, 
        NET_CC_CONFIG47, NET_CC_CONFIG48, NET_CC_CONFIG49, 
        NET_CC_CONFIG50, NET_CC_CONFIG51, NET_CC_CONFIG52, 
        NET_CC_CONFIG53, NET_CC_CONFIG54, NET_CC_CONFIG55, 
        NET_CC_CONFIG56, NET_CC_CONFIG57, NET_CC_CONFIG58, 
        NET_CC_CONFIG59, NET_CC_CONFIG60, NET_CC_CONFIG61, 
        NET_CC_CONFIG62, NET_CC_CONFIG63, NET_CC_CONFIG64, 
        NET_CC_CONFIG65, NET_CC_CONFIG66, NET_CC_CONFIG67, 
        NET_CC_CONFIG68, NET_CC_CONFIG69, NET_CC_CONFIG70, 
        NET_CC_CONFIG71, NET_CC_CONFIG72, NET_CC_CONFIG73, 
        NET_CC_CONFIG74, NET_CC_CONFIG75, NET_CC_CONFIG76, 
        NET_CC_CONFIG77, NET_CC_CONFIG78, NET_CC_CONFIG79, 
        NET_CC_CONFIG80, NET_CC_CONFIG81, NET_CC_CONFIG82, 
        NET_CC_CONFIG83, NET_CC_CONFIG84, NET_CC_CONFIG85, 
        NET_CC_CONFIG86, NET_CC_CONFIG87, NET_CC_CONFIG88, 
        NET_CC_CONFIG89, NET_CC_CONFIG90, NET_CC_CONFIG91, 
        NET_CC_CONFIG92, NET_CC_CONFIG93, NET_CC_CONFIG94, 
        NET_CC_CONFIG95, NET_CC_CONFIG96, NET_CC_CONFIG97, 
        NET_CC_CONFIG98, NET_CC_CONFIG99, CI_TO_CO100, 
        CI_TO_CO101, NET_CC_CONFIG102, NET_CC_CONFIG103, 
        NET_CC_CONFIG104, NET_CC_CONFIG105, NET_CC_CONFIG106, 
        NET_CC_CONFIG107, NET_CC_CONFIG108, NET_CC_CONFIG109, 
        NET_CC_CONFIG110, NET_CC_CONFIG111, NET_CC_CONFIG112, 
        NET_CC_CONFIG113, NET_CC_CONFIG114, NET_CC_CONFIG115, 
        NET_CC_CONFIG116, NET_CC_CONFIG117, NET_CC_CONFIG118, 
        NET_CC_CONFIG119, NET_CC_CONFIG120, NET_CC_CONFIG121, 
        NET_CC_CONFIG122, NET_CC_CONFIG123, NET_CC_CONFIG124, 
        NET_CC_CONFIG125, NET_CC_CONFIG126, NET_CC_CONFIG127, 
        NET_CC_CONFIG128, NET_CC_CONFIG129, NET_CC_CONFIG130, 
        NET_CC_CONFIG131, NET_CC_CONFIG132, NET_CC_CONFIG133, 
        NET_CC_CONFIG134, NET_CC_CONFIG135, NET_CC_CONFIG136, 
        NET_CC_CONFIG137, NET_CC_CONFIG138, NET_CC_CONFIG139, 
        NET_CC_CONFIG140, NET_CC_CONFIG141, NET_CC_CONFIG142, 
        NET_CC_CONFIG143, NET_CC_CONFIG144, NET_CC_CONFIG145, 
        NET_CC_CONFIG146, NET_CC_CONFIG147, NET_CC_CONFIG148, 
        NET_CC_CONFIG149, NET_CC_CONFIG150, NET_CC_CONFIG151, 
        NET_CC_CONFIG152, NET_CC_CONFIG153, NET_CC_CONFIG154, 
        NET_CC_CONFIG155, NET_CC_CONFIG156, NET_CC_CONFIG157, 
        NET_CC_CONFIG158, NET_CC_CONFIG159, NET_CC_CONFIG160, 
        NET_CC_CONFIG161, NET_CC_CONFIG162, NET_CC_CONFIG163, 
        NET_CC_CONFIG164, NET_CC_CONFIG165, NET_CC_CONFIG166, 
        NET_CC_CONFIG167, NET_CC_CONFIG168, NET_CC_CONFIG169, 
        NET_CC_CONFIG170, NET_CC_CONFIG171, NET_CC_CONFIG172, 
        NET_CC_CONFIG173, NET_CC_CONFIG174, NET_CC_CONFIG175, 
        NET_CC_CONFIG176, NET_CC_CONFIG177, NET_CC_CONFIG178, 
        NET_CC_CONFIG179, NET_CC_CONFIG180, NET_CC_CONFIG181, 
        NET_CC_CONFIG182, NET_CC_CONFIG183, NET_CC_CONFIG184, 
        NET_CC_CONFIG185, NET_CC_CONFIG186, NET_CC_CONFIG187, 
        NET_CC_CONFIG188, NET_CC_CONFIG189, NET_CC_CONFIG190, 
        NET_CC_CONFIG191, NET_CC_CONFIG192, NET_CC_CONFIG193, 
        NET_CC_CONFIG194, CI_TO_CO195, CI_TO_CO196, 
        NET_CC_CONFIG197, NET_CC_CONFIG198, NET_CC_CONFIG199, 
        NET_CC_CONFIG200, NET_CC_CONFIG201, NET_CC_CONFIG202, 
        NET_CC_CONFIG203, NET_CC_CONFIG204, NET_CC_CONFIG205, 
        NET_CC_CONFIG206, NET_CC_CONFIG207, NET_CC_CONFIG208, 
        NET_CC_CONFIG209, NET_CC_CONFIG210, NET_CC_CONFIG211, 
        NET_CC_CONFIG212, NET_CC_CONFIG213, NET_CC_CONFIG214, 
        NET_CC_CONFIG215, NET_CC_CONFIG216, NET_CC_CONFIG217, 
        NET_CC_CONFIG218, NET_CC_CONFIG219, NET_CC_CONFIG220, 
        NET_CC_CONFIG221, NET_CC_CONFIG222, NET_CC_CONFIG223, 
        NET_CC_CONFIG224, NET_CC_CONFIG225, NET_CC_CONFIG226, 
        NET_CC_CONFIG227, NET_CC_CONFIG228, NET_CC_CONFIG229, 
        NET_CC_CONFIG230, NET_CC_CONFIG231, NET_CC_CONFIG232, 
        NET_CC_CONFIG233, NET_CC_CONFIG234, NET_CC_CONFIG235, 
        NET_CC_CONFIG236, NET_CC_CONFIG237, NET_CC_CONFIG238, 
        NET_CC_CONFIG239, NET_CC_CONFIG240, NET_CC_CONFIG241, 
        NET_CC_CONFIG242, NET_CC_CONFIG243, NET_CC_CONFIG244, 
        NET_CC_CONFIG245, NET_CC_CONFIG246, NET_CC_CONFIG247, 
        NET_CC_CONFIG248, NET_CC_CONFIG249, NET_CC_CONFIG250, 
        NET_CC_CONFIG251, NET_CC_CONFIG252, NET_CC_CONFIG253, 
        NET_CC_CONFIG254, NET_CC_CONFIG255, NET_CC_CONFIG256, 
        NET_CC_CONFIG257, NET_CC_CONFIG258, NET_CC_CONFIG259, 
        NET_CC_CONFIG260, NET_CC_CONFIG261, NET_CC_CONFIG262, 
        NET_CC_CONFIG263, NET_CC_CONFIG264, NET_CC_CONFIG265, 
        NET_CC_CONFIG266, NET_CC_CONFIG267, NET_CC_CONFIG268, 
        NET_CC_CONFIG269, NET_CC_CONFIG270, NET_CC_CONFIG271, 
        NET_CC_CONFIG272, NET_CC_CONFIG273, NET_CC_CONFIG274, 
        NET_CC_CONFIG275, NET_CC_CONFIG276, NET_CC_CONFIG277, 
        NET_CC_CONFIG278, NET_CC_CONFIG279, NET_CC_CONFIG280, 
        NET_CC_CONFIG281, NET_CC_CONFIG282, NET_CC_CONFIG283, 
        NET_CC_CONFIG284, NET_CC_CONFIG285, NET_CC_CONFIG286, 
        NET_CC_CONFIG287, NET_CC_CONFIG288, NET_CC_CONFIG289, 
        NET_CC_CONFIG290, NET_CC_CONFIG291, NET_CC_CONFIG292, 
        CI_TO_CO293, CI_TO_CO294, NET_CC_CONFIG295, 
        NET_CC_CONFIG296, NET_CC_CONFIG297, NET_CC_CONFIG298, 
        NET_CC_CONFIG299, NET_CC_CONFIG300, NET_CC_CONFIG301, 
        NET_CC_CONFIG302, NET_CC_CONFIG303, NET_CC_CONFIG304, 
        NET_CC_CONFIG305, NET_CC_CONFIG306, NET_CC_CONFIG307, 
        NET_CC_CONFIG308, NET_CC_CONFIG309, NET_CC_CONFIG310, 
        NET_CC_CONFIG311, NET_CC_CONFIG312, NET_CC_CONFIG313, 
        NET_CC_CONFIG314, NET_CC_CONFIG315, NET_CC_CONFIG316, 
        NET_CC_CONFIG317, NET_CC_CONFIG318, NET_CC_CONFIG319, 
        NET_CC_CONFIG320, NET_CC_CONFIG321, NET_CC_CONFIG322, 
        NET_CC_CONFIG323, NET_CC_CONFIG324, NET_CC_CONFIG325, 
        NET_CC_CONFIG326, NET_CC_CONFIG327, NET_CC_CONFIG328, 
        NET_CC_CONFIG329, NET_CC_CONFIG330, NET_CC_CONFIG331, 
        NET_CC_CONFIG332, NET_CC_CONFIG333, NET_CC_CONFIG334, 
        NET_CC_CONFIG335, NET_CC_CONFIG336, NET_CC_CONFIG337, 
        NET_CC_CONFIG338, NET_CC_CONFIG339, NET_CC_CONFIG340, 
        NET_CC_CONFIG341, NET_CC_CONFIG342, NET_CC_CONFIG343, 
        NET_CC_CONFIG344, NET_CC_CONFIG345, NET_CC_CONFIG346, 
        NET_CC_CONFIG347, NET_CC_CONFIG348, NET_CC_CONFIG349, 
        NET_CC_CONFIG350, NET_CC_CONFIG351, NET_CC_CONFIG352, 
        NET_CC_CONFIG353, NET_CC_CONFIG354, NET_CC_CONFIG355, 
        NET_CC_CONFIG356, NET_CC_CONFIG357, NET_CC_CONFIG358, 
        NET_CC_CONFIG359, NET_CC_CONFIG360, NET_CC_CONFIG361, 
        NET_CC_CONFIG362, NET_CC_CONFIG363, NET_CC_CONFIG364, 
        NET_CC_CONFIG365, NET_CC_CONFIG366, NET_CC_CONFIG367, 
        NET_CC_CONFIG368, NET_CC_CONFIG369, NET_CC_CONFIG370, 
        NET_CC_CONFIG371, NET_CC_CONFIG372, NET_CC_CONFIG373, 
        NET_CC_CONFIG374, NET_CC_CONFIG375, NET_CC_CONFIG376, 
        NET_CC_CONFIG377, NET_CC_CONFIG378, NET_CC_CONFIG379, 
        NET_CC_CONFIG380, NET_CC_CONFIG381, NET_CC_CONFIG382, 
        NET_CC_CONFIG383, NET_CC_CONFIG384, NET_CC_CONFIG385, 
        NET_CC_CONFIG386, NET_CC_CONFIG387, NET_CC_CONFIG388, 
        NET_CC_CONFIG389, NET_CC_CONFIG390, CI_TO_CO391, 
        CI_TO_CO392, NET_CC_CONFIG393, NET_CC_CONFIG394, 
        NET_CC_CONFIG395, NET_CC_CONFIG396, NET_CC_CONFIG397, 
        NET_CC_CONFIG398, NET_CC_CONFIG399, NET_CC_CONFIG400, 
        NET_CC_CONFIG401, NET_CC_CONFIG402, NET_CC_CONFIG403, 
        NET_CC_CONFIG404, NET_CC_CONFIG405, NET_CC_CONFIG406, 
        NET_CC_CONFIG407, NET_CC_CONFIG408, NET_CC_CONFIG409, 
        NET_CC_CONFIG410, NET_CC_CONFIG411, NET_CC_CONFIG412, 
        NET_CC_CONFIG413, NET_CC_CONFIG414, NET_CC_CONFIG415, 
        NET_CC_CONFIG416, NET_CC_CONFIG417, NET_CC_CONFIG418, 
        NET_CC_CONFIG419, NET_CC_CONFIG420, NET_CC_CONFIG421, 
        NET_CC_CONFIG422, NET_CC_CONFIG423, NET_CC_CONFIG424, 
        NET_CC_CONFIG425, NET_CC_CONFIG426, NET_CC_CONFIG427, 
        NET_CC_CONFIG428, NET_CC_CONFIG429, NET_CC_CONFIG430, 
        NET_CC_CONFIG431, NET_CC_CONFIG432, NET_CC_CONFIG433, 
        NET_CC_CONFIG434, NET_CC_CONFIG435, NET_CC_CONFIG436, 
        NET_CC_CONFIG437, NET_CC_CONFIG438, NET_CC_CONFIG439, 
        NET_CC_CONFIG440, NET_CC_CONFIG441, NET_CC_CONFIG442, 
        NET_CC_CONFIG443, NET_CC_CONFIG444, NET_CC_CONFIG445, 
        NET_CC_CONFIG446, NET_CC_CONFIG447, NET_CC_CONFIG448, 
        NET_CC_CONFIG449, NET_CC_CONFIG450, NET_CC_CONFIG451, 
        NET_CC_CONFIG452, NET_CC_CONFIG453, NET_CC_CONFIG454, 
        NET_CC_CONFIG455, NET_CC_CONFIG456, NET_CC_CONFIG457, 
        NET_CC_CONFIG458, NET_CC_CONFIG459, NET_CC_CONFIG460, 
        NET_CC_CONFIG461, NET_CC_CONFIG462, NET_CC_CONFIG463, 
        NET_CC_CONFIG464, NET_CC_CONFIG465, NET_CC_CONFIG466, 
        NET_CC_CONFIG467, NET_CC_CONFIG468, NET_CC_CONFIG469, 
        NET_CC_CONFIG470, NET_CC_CONFIG471, NET_CC_CONFIG472, 
        NET_CC_CONFIG473, NET_CC_CONFIG474, NET_CC_CONFIG475, 
        NET_CC_CONFIG476, CI_TO_CO477, NET_CC_CONFIG478, 
        NET_CC_CONFIG479, NET_CC_CONFIG480, NET_CC_CONFIG481, 
        NET_CC_CONFIG482, NET_CC_CONFIG483, NET_CC_CONFIG484, 
        NET_CC_CONFIG485, NET_CC_CONFIG486, NET_CC_CONFIG487, 
        NET_CC_CONFIG488, NET_CC_CONFIG489, NET_CC_CONFIG490, 
        NET_CC_CONFIG491, NET_CC_CONFIG492, NET_CC_CONFIG493, 
        NET_CC_CONFIG494, NET_CC_CONFIG495, NET_CC_CONFIG496, 
        NET_CC_CONFIG497, NET_CC_CONFIG498, NET_CC_CONFIG499, 
        NET_CC_CONFIG500, NET_CC_CONFIG501, NET_CC_CONFIG502, 
        NET_CC_CONFIG503, NET_CC_CONFIG504, NET_CC_CONFIG505, 
        NET_CC_CONFIG506, NET_CC_CONFIG507, NET_CC_CONFIG508, 
        NET_CC_CONFIG509, NET_CC_CONFIG510, NET_CC_CONFIG511, 
        NET_CC_CONFIG512, NET_CC_CONFIG513, NET_CC_CONFIG514, 
        NET_CC_CONFIG515, NET_CC_CONFIG516, NET_CC_CONFIG517, 
        NET_CC_CONFIG518, NET_CC_CONFIG519, NET_CC_CONFIG520, 
        NET_CC_CONFIG521, NET_CC_CONFIG522, NET_CC_CONFIG523, 
        NET_CC_CONFIG524, NET_CC_CONFIG525, NET_CC_CONFIG526, 
        NET_CC_CONFIG527, NET_CC_CONFIG528, NET_CC_CONFIG529, 
        NET_CC_CONFIG530, NET_CC_CONFIG531, NET_CC_CONFIG532, 
        NET_CC_CONFIG533, NET_CC_CONFIG534, CI_TO_CO535, 
        NET_CC_CONFIG536, NET_CC_CONFIG537, NET_CC_CONFIG538, 
        NET_CC_CONFIG539, NET_CC_CONFIG540, NET_CC_CONFIG541, 
        NET_CC_CONFIG542, NET_CC_CONFIG543, NET_CC_CONFIG544, 
        NET_CC_CONFIG545, NET_CC_CONFIG546, NET_CC_CONFIG547, 
        NET_CC_CONFIG548, NET_CC_CONFIG549, NET_CC_CONFIG550, 
        NET_CC_CONFIG551, NET_CC_CONFIG552, NET_CC_CONFIG553, 
        NET_CC_CONFIG554, NET_CC_CONFIG555, NET_CC_CONFIG556, 
        NET_CC_CONFIG557, NET_CC_CONFIG558, NET_CC_CONFIG559, 
        NET_CC_CONFIG560, NET_CC_CONFIG561, NET_CC_CONFIG562, 
        NET_CC_CONFIG563, NET_CC_CONFIG564, NET_CC_CONFIG565, 
        NET_CC_CONFIG566, NET_CC_CONFIG567, NET_CC_CONFIG568, 
        NET_CC_CONFIG569, NET_CC_CONFIG570, NET_CC_CONFIG571, 
        NET_CC_CONFIG572, NET_CC_CONFIG573, NET_CC_CONFIG574, 
        NET_CC_CONFIG575, NET_CC_CONFIG576, NET_CC_CONFIG577, 
        NET_CC_CONFIG578, NET_CC_CONFIG579, NET_CC_CONFIG580, 
        NET_CC_CONFIG581, NET_CC_CONFIG582, NET_CC_CONFIG583, 
        NET_CC_CONFIG584, NET_CC_CONFIG585, NET_CC_CONFIG586, 
        NET_CC_CONFIG587, NET_CC_CONFIG588, NET_CC_CONFIG589, 
        NET_CC_CONFIG590, NET_CC_CONFIG591, NET_CC_CONFIG592, 
        NET_CC_CONFIG593, NET_CC_CONFIG594, NET_CC_CONFIG595, 
        NET_CC_CONFIG596, NET_CC_CONFIG597, NET_CC_CONFIG598, 
        NET_CC_CONFIG599, NET_CC_CONFIG600, NET_CC_CONFIG601, 
        NET_CC_CONFIG602, NET_CC_CONFIG603, NET_CC_CONFIG604, 
        NET_CC_CONFIG605, NET_CC_CONFIG606, NET_CC_CONFIG607, 
        NET_CC_CONFIG608, NET_CC_CONFIG609, NET_CC_CONFIG610, 
        NET_CC_CONFIG611, NET_CC_CONFIG612, NET_CC_CONFIG613, 
        NET_CC_CONFIG614, NET_CC_CONFIG615, NET_CC_CONFIG616, 
        NET_CC_CONFIG617, NET_CC_CONFIG618, NET_CC_CONFIG619, 
        NET_CC_CONFIG620, NET_CC_CONFIG621, NET_CC_CONFIG622, 
        CI_TO_CO623, CI_TO_CO624, NET_CC_CONFIG625, 
        NET_CC_CONFIG626, NET_CC_CONFIG627, NET_CC_CONFIG628, 
        NET_CC_CONFIG629, NET_CC_CONFIG630, NET_CC_CONFIG631, 
        NET_CC_CONFIG632, NET_CC_CONFIG633, NET_CC_CONFIG634, 
        NET_CC_CONFIG635, NET_CC_CONFIG636, NET_CC_CONFIG637, 
        NET_CC_CONFIG638, NET_CC_CONFIG639, NET_CC_CONFIG640, 
        NET_CC_CONFIG641, NET_CC_CONFIG642, NET_CC_CONFIG643, 
        NET_CC_CONFIG644, NET_CC_CONFIG645, NET_CC_CONFIG646, 
        NET_CC_CONFIG647, NET_CC_CONFIG648, NET_CC_CONFIG649, 
        NET_CC_CONFIG650, NET_CC_CONFIG651, NET_CC_CONFIG652, 
        NET_CC_CONFIG653, NET_CC_CONFIG654, NET_CC_CONFIG655, 
        NET_CC_CONFIG656, NET_CC_CONFIG657, NET_CC_CONFIG658, 
        NET_CC_CONFIG659, NET_CC_CONFIG660, NET_CC_CONFIG661, 
        NET_CC_CONFIG662, NET_CC_CONFIG663, NET_CC_CONFIG664, 
        NET_CC_CONFIG665, NET_CC_CONFIG666, NET_CC_CONFIG667, 
        NET_CC_CONFIG668, NET_CC_CONFIG669, NET_CC_CONFIG670, 
        NET_CC_CONFIG671, NET_CC_CONFIG672, NET_CC_CONFIG673, 
        NET_CC_CONFIG674, NET_CC_CONFIG675, NET_CC_CONFIG676, 
        NET_CC_CONFIG677, NET_CC_CONFIG678, NET_CC_CONFIG679, 
        NET_CC_CONFIG680, NET_CC_CONFIG681, NET_CC_CONFIG682, 
        NET_CC_CONFIG683, NET_CC_CONFIG684, NET_CC_CONFIG685, 
        NET_CC_CONFIG686, NET_CC_CONFIG687, NET_CC_CONFIG688, 
        NET_CC_CONFIG689, NET_CC_CONFIG690, NET_CC_CONFIG691, 
        NET_CC_CONFIG692, NET_CC_CONFIG693, NET_CC_CONFIG694, 
        NET_CC_CONFIG695, NET_CC_CONFIG696, NET_CC_CONFIG697, 
        NET_CC_CONFIG698, NET_CC_CONFIG699, NET_CC_CONFIG700, 
        NET_CC_CONFIG701, NET_CC_CONFIG702, NET_CC_CONFIG703, 
        NET_CC_CONFIG704, NET_CC_CONFIG705, NET_CC_CONFIG706, 
        NET_CC_CONFIG707, NET_CC_CONFIG708, NET_CC_CONFIG709, 
        NET_CC_CONFIG710, NET_CC_CONFIG711, NET_CC_CONFIG712, 
        NET_CC_CONFIG713, NET_CC_CONFIG714, NET_CC_CONFIG715, 
        NET_CC_CONFIG716, NET_CC_CONFIG717, NET_CC_CONFIG718, 
        NET_CC_CONFIG719, NET_CC_CONFIG720, CI_TO_CO721, 
        CI_TO_CO722, NET_CC_CONFIG723, NET_CC_CONFIG724, 
        NET_CC_CONFIG725, NET_CC_CONFIG726, NET_CC_CONFIG727, 
        NET_CC_CONFIG728, NET_CC_CONFIG729, NET_CC_CONFIG730, 
        NET_CC_CONFIG731, NET_CC_CONFIG732, NET_CC_CONFIG733, 
        NET_CC_CONFIG734, NET_CC_CONFIG735, NET_CC_CONFIG736, 
        NET_CC_CONFIG737, NET_CC_CONFIG738, NET_CC_CONFIG739, 
        NET_CC_CONFIG740, NET_CC_CONFIG741, NET_CC_CONFIG742, 
        NET_CC_CONFIG743, NET_CC_CONFIG744, NET_CC_CONFIG745, 
        NET_CC_CONFIG746, NET_CC_CONFIG747, NET_CC_CONFIG748, 
        NET_CC_CONFIG749, NET_CC_CONFIG750, NET_CC_CONFIG751, 
        NET_CC_CONFIG752, NET_CC_CONFIG753, NET_CC_CONFIG754, 
        NET_CC_CONFIG755, NET_CC_CONFIG756, NET_CC_CONFIG757, 
        NET_CC_CONFIG758, NET_CC_CONFIG759, NET_CC_CONFIG760, 
        NET_CC_CONFIG761, NET_CC_CONFIG762, NET_CC_CONFIG763, 
        NET_CC_CONFIG764, NET_CC_CONFIG765, NET_CC_CONFIG766, 
        NET_CC_CONFIG767, NET_CC_CONFIG768, NET_CC_CONFIG769, 
        NET_CC_CONFIG770, NET_CC_CONFIG771, NET_CC_CONFIG772, 
        NET_CC_CONFIG773, NET_CC_CONFIG774, NET_CC_CONFIG775, 
        NET_CC_CONFIG776, NET_CC_CONFIG777, NET_CC_CONFIG778, 
        NET_CC_CONFIG779, NET_CC_CONFIG780, NET_CC_CONFIG781, 
        NET_CC_CONFIG782, NET_CC_CONFIG783, NET_CC_CONFIG784, 
        NET_CC_CONFIG785, NET_CC_CONFIG786, NET_CC_CONFIG787, 
        NET_CC_CONFIG788, NET_CC_CONFIG789, NET_CC_CONFIG790, 
        NET_CC_CONFIG791, NET_CC_CONFIG792, NET_CC_CONFIG793, 
        NET_CC_CONFIG794, NET_CC_CONFIG795, NET_CC_CONFIG796, 
        NET_CC_CONFIG797, NET_CC_CONFIG798, NET_CC_CONFIG799, 
        NET_CC_CONFIG800, NET_CC_CONFIG801, NET_CC_CONFIG802, 
        NET_CC_CONFIG803, NET_CC_CONFIG804, NET_CC_CONFIG805, 
        NET_CC_CONFIG806, NET_CC_CONFIG807, NET_CC_CONFIG808, 
        NET_CC_CONFIG809, NET_CC_CONFIG810, NET_CC_CONFIG811, 
        NET_CC_CONFIG812, NET_CC_CONFIG813, NET_CC_CONFIG814, 
        NET_CC_CONFIG815, NET_CC_CONFIG816, NET_CC_CONFIG817, 
        NET_CC_CONFIG818, CI_TO_CO819, CI_TO_CO820, 
        NET_CC_CONFIG821, NET_CC_CONFIG822, NET_CC_CONFIG823, 
        NET_CC_CONFIG824, NET_CC_CONFIG825, NET_CC_CONFIG826, 
        NET_CC_CONFIG827, NET_CC_CONFIG828, NET_CC_CONFIG829, 
        NET_CC_CONFIG830, NET_CC_CONFIG831, NET_CC_CONFIG832, 
        NET_CC_CONFIG833, NET_CC_CONFIG834, NET_CC_CONFIG835, 
        NET_CC_CONFIG836, NET_CC_CONFIG837, NET_CC_CONFIG838, 
        NET_CC_CONFIG839, NET_CC_CONFIG840, NET_CC_CONFIG841, 
        NET_CC_CONFIG842, NET_CC_CONFIG843, NET_CC_CONFIG844, 
        NET_CC_CONFIG845, NET_CC_CONFIG846, NET_CC_CONFIG847, 
        NET_CC_CONFIG848, NET_CC_CONFIG849, NET_CC_CONFIG850, 
        NET_CC_CONFIG851, NET_CC_CONFIG852, NET_CC_CONFIG853, 
        NET_CC_CONFIG854, NET_CC_CONFIG855, NET_CC_CONFIG856, 
        NET_CC_CONFIG857, NET_CC_CONFIG858, NET_CC_CONFIG859, 
        NET_CC_CONFIG860, NET_CC_CONFIG861, NET_CC_CONFIG862, 
        NET_CC_CONFIG863, NET_CC_CONFIG864, NET_CC_CONFIG865, 
        NET_CC_CONFIG866, NET_CC_CONFIG867, NET_CC_CONFIG868, 
        NET_CC_CONFIG869, NET_CC_CONFIG870, NET_CC_CONFIG871, 
        NET_CC_CONFIG872, NET_CC_CONFIG873, NET_CC_CONFIG874, 
        NET_CC_CONFIG875, NET_CC_CONFIG876, NET_CC_CONFIG877, 
        NET_CC_CONFIG878, NET_CC_CONFIG879, NET_CC_CONFIG880, 
        NET_CC_CONFIG881, NET_CC_CONFIG882, NET_CC_CONFIG883, 
        NET_CC_CONFIG884, NET_CC_CONFIG885, NET_CC_CONFIG886, 
        NET_CC_CONFIG887, NET_CC_CONFIG888, NET_CC_CONFIG889, 
        NET_CC_CONFIG890, NET_CC_CONFIG891, NET_CC_CONFIG892, 
        NET_CC_CONFIG893, NET_CC_CONFIG894, NET_CC_CONFIG895, 
        NET_CC_CONFIG896, NET_CC_CONFIG897, NET_CC_CONFIG898, 
        NET_CC_CONFIG899, NET_CC_CONFIG900, NET_CC_CONFIG901, 
        NET_CC_CONFIG902, NET_CC_CONFIG903, NET_CC_CONFIG904, 
        NET_CC_CONFIG905, NET_CC_CONFIG906, NET_CC_CONFIG907, 
        NET_CC_CONFIG908, NET_CC_CONFIG909, NET_CC_CONFIG910, 
        NET_CC_CONFIG911, NET_CC_CONFIG912, NET_CC_CONFIG913, 
        NET_CC_CONFIG914, NET_CC_CONFIG915, NET_CC_CONFIG916, 
        NET_CC_CONFIG917, NET_CC_CONFIG918, NET_CC_CONFIG919, 
        CI_TO_CO920, CI_TO_CO921, CI_TO_CO922, NET_CC_CONFIG923, 
        NET_CC_CONFIG924, NET_CC_CONFIG925, NET_CC_CONFIG926, 
        NET_CC_CONFIG927, NET_CC_CONFIG928, NET_CC_CONFIG929, 
        NET_CC_CONFIG930, NET_CC_CONFIG931, NET_CC_CONFIG932, 
        NET_CC_CONFIG933, NET_CC_CONFIG934, NET_CC_CONFIG935, 
        NET_CC_CONFIG936, NET_CC_CONFIG937, NET_CC_CONFIG938, 
        NET_CC_CONFIG939, NET_CC_CONFIG940, NET_CC_CONFIG941, 
        NET_CC_CONFIG942, NET_CC_CONFIG943, NET_CC_CONFIG944, 
        NET_CC_CONFIG945, NET_CC_CONFIG946, NET_CC_CONFIG947, 
        NET_CC_CONFIG948, NET_CC_CONFIG949, NET_CC_CONFIG950, 
        NET_CC_CONFIG951, NET_CC_CONFIG952, NET_CC_CONFIG953, 
        NET_CC_CONFIG954, NET_CC_CONFIG955, NET_CC_CONFIG956, 
        NET_CC_CONFIG957, NET_CC_CONFIG958, NET_CC_CONFIG959, 
        NET_CC_CONFIG960, NET_CC_CONFIG961, NET_CC_CONFIG962, 
        NET_CC_CONFIG963, NET_CC_CONFIG964, NET_CC_CONFIG965, 
        NET_CC_CONFIG966, NET_CC_CONFIG967, NET_CC_CONFIG968, 
        NET_CC_CONFIG969, NET_CC_CONFIG970, NET_CC_CONFIG971, 
        NET_CC_CONFIG972, NET_CC_CONFIG973, NET_CC_CONFIG974, 
        NET_CC_CONFIG975, NET_CC_CONFIG976, NET_CC_CONFIG977, 
        NET_CC_CONFIG978, NET_CC_CONFIG979, NET_CC_CONFIG980, 
        NET_CC_CONFIG981, NET_CC_CONFIG982, NET_CC_CONFIG983, 
        NET_CC_CONFIG984, NET_CC_CONFIG985, NET_CC_CONFIG986, 
        NET_CC_CONFIG987, NET_CC_CONFIG988, NET_CC_CONFIG989, 
        NET_CC_CONFIG990, NET_CC_CONFIG991, NET_CC_CONFIG992, 
        NET_CC_CONFIG993, NET_CC_CONFIG994, NET_CC_CONFIG995, 
        NET_CC_CONFIG996, NET_CC_CONFIG997, NET_CC_CONFIG998, 
        NET_CC_CONFIG999, NET_CC_CONFIG1000, NET_CC_CONFIG1001, 
        NET_CC_CONFIG1002, NET_CC_CONFIG1003, NET_CC_CONFIG1004, 
        NET_CC_CONFIG1005, NET_CC_CONFIG1006, NET_CC_CONFIG1007, 
        NET_CC_CONFIG1008, NET_CC_CONFIG1009, NET_CC_CONFIG1010, 
        NET_CC_CONFIG1011, NET_CC_CONFIG1012, NET_CC_CONFIG1013, 
        NET_CC_CONFIG1014, NET_CC_CONFIG1015, NET_CC_CONFIG1016, 
        NET_CC_CONFIG1017, NET_CC_CONFIG1018, CI_TO_CO1019, 
        CI_TO_CO1020, NET_CC_CONFIG1021, NET_CC_CONFIG1022, 
        NET_CC_CONFIG1023, NET_CC_CONFIG1024, NET_CC_CONFIG1025, 
        NET_CC_CONFIG1026, NET_CC_CONFIG1027, NET_CC_CONFIG1028, 
        NET_CC_CONFIG1029, NET_CC_CONFIG1030, NET_CC_CONFIG1031, 
        NET_CC_CONFIG1032, NET_CC_CONFIG1033, NET_CC_CONFIG1034, 
        NET_CC_CONFIG1035, NET_CC_CONFIG1036, NET_CC_CONFIG1037, 
        NET_CC_CONFIG1038, NET_CC_CONFIG1039, NET_CC_CONFIG1040, 
        NET_CC_CONFIG1041, NET_CC_CONFIG1042, NET_CC_CONFIG1043, 
        NET_CC_CONFIG1044, NET_CC_CONFIG1045, NET_CC_CONFIG1046, 
        NET_CC_CONFIG1047, NET_CC_CONFIG1048, NET_CC_CONFIG1049, 
        NET_CC_CONFIG1050, NET_CC_CONFIG1051, NET_CC_CONFIG1052, 
        NET_CC_CONFIG1053, NET_CC_CONFIG1054, NET_CC_CONFIG1055, 
        NET_CC_CONFIG1056, NET_CC_CONFIG1057, NET_CC_CONFIG1058, 
        NET_CC_CONFIG1059, NET_CC_CONFIG1060, NET_CC_CONFIG1061, 
        NET_CC_CONFIG1062, NET_CC_CONFIG1063, NET_CC_CONFIG1064, 
        NET_CC_CONFIG1065, NET_CC_CONFIG1066, NET_CC_CONFIG1067, 
        NET_CC_CONFIG1068, NET_CC_CONFIG1069, NET_CC_CONFIG1070, 
        NET_CC_CONFIG1071, NET_CC_CONFIG1072, NET_CC_CONFIG1073, 
        NET_CC_CONFIG1074, NET_CC_CONFIG1075, NET_CC_CONFIG1076, 
        NET_CC_CONFIG1077, NET_CC_CONFIG1078, NET_CC_CONFIG1079, 
        NET_CC_CONFIG1080, NET_CC_CONFIG1081, NET_CC_CONFIG1082, 
        NET_CC_CONFIG1083, NET_CC_CONFIG1084, NET_CC_CONFIG1085, 
        NET_CC_CONFIG1086, NET_CC_CONFIG1087, NET_CC_CONFIG1088, 
        NET_CC_CONFIG1089, NET_CC_CONFIG1090, NET_CC_CONFIG1091, 
        NET_CC_CONFIG1092, NET_CC_CONFIG1093, NET_CC_CONFIG1094, 
        NET_CC_CONFIG1095, NET_CC_CONFIG1096, NET_CC_CONFIG1097, 
        NET_CC_CONFIG1098, NET_CC_CONFIG1099, NET_CC_CONFIG1100, 
        NET_CC_CONFIG1101, NET_CC_CONFIG1102, NET_CC_CONFIG1103, 
        NET_CC_CONFIG1104, NET_CC_CONFIG1105, NET_CC_CONFIG1106, 
        NET_CC_CONFIG1107, NET_CC_CONFIG1108, NET_CC_CONFIG1109, 
        NET_CC_CONFIG1110, NET_CC_CONFIG1111, NET_CC_CONFIG1112, 
        NET_CC_CONFIG1113, CI_TO_CO1114, NET_CC_CONFIG1115, 
        NET_CC_CONFIG1116, NET_CC_CONFIG1117, NET_CC_CONFIG1118, 
        NET_CC_CONFIG1119, NET_CC_CONFIG1120, NET_CC_CONFIG1121, 
        NET_CC_CONFIG1122, NET_CC_CONFIG1123, NET_CC_CONFIG1124, 
        NET_CC_CONFIG1125, NET_CC_CONFIG1126, NET_CC_CONFIG1127, 
        NET_CC_CONFIG1128, NET_CC_CONFIG1129, NET_CC_CONFIG1130, 
        NET_CC_CONFIG1131, NET_CC_CONFIG1132, NET_CC_CONFIG1133, 
        NET_CC_CONFIG1134, NET_CC_CONFIG1135, NET_CC_CONFIG1136, 
        NET_CC_CONFIG1137, NET_CC_CONFIG1138, NET_CC_CONFIG1139, 
        NET_CC_CONFIG1140, NET_CC_CONFIG1141, NET_CC_CONFIG1142, 
        NET_CC_CONFIG1143, NET_CC_CONFIG1144, NET_CC_CONFIG1145, 
        NET_CC_CONFIG1146, NET_CC_CONFIG1147, NET_CC_CONFIG1148, 
        NET_CC_CONFIG1149, NET_CC_CONFIG1150, NET_CC_CONFIG1151, 
        NET_CC_CONFIG1152, NET_CC_CONFIG1153, NET_CC_CONFIG1154, 
        NET_CC_CONFIG1155, NET_CC_CONFIG1156, NET_CC_CONFIG1157, 
        NET_CC_CONFIG1158, NET_CC_CONFIG1159, NET_CC_CONFIG1160, 
        NET_CC_CONFIG1161, NET_CC_CONFIG1162, NET_CC_CONFIG1163, 
        NET_CC_CONFIG1164, NET_CC_CONFIG1165, AFLSDF_VCC, 
        AFLSDF_GND, \AFLSDF_INV_0\, \AFLSDF_INV_1\, 
        \AFLSDF_INV_2\, \AFLSDF_INV_3\, \AFLSDF_INV_4\, 
        \AFLSDF_INV_5\, \AFLSDF_INV_6\, \AFLSDF_INV_7\, 
        \AFLSDF_INV_8\, \AFLSDF_INV_9\, \AFLSDF_INV_10\, 
        \AFLSDF_INV_11\, \AFLSDF_INV_12\, \AFLSDF_INV_13\, 
        \AFLSDF_INV_14\, \AFLSDF_INV_15\, \AFLSDF_INV_16\, 
        \AFLSDF_INV_17\, \AFLSDF_INV_18\, \AFLSDF_INV_19\, 
        \AFLSDF_INV_20\, \AFLSDF_INV_21\, \AFLSDF_INV_22\, 
        \AFLSDF_INV_23\, \AFLSDF_INV_24\, \AFLSDF_INV_25\, 
        \AFLSDF_INV_26\, \AFLSDF_INV_27\, \AFLSDF_INV_28\, 
        \AFLSDF_INV_29\, \AFLSDF_INV_30\, \AFLSDF_INV_31\, 
        \AFLSDF_INV_32\, \AFLSDF_INV_33\, \AFLSDF_INV_34\, 
        \AFLSDF_INV_35\, \AFLSDF_INV_36\, \AFLSDF_INV_37\, 
        \AFLSDF_INV_38\, \AFLSDF_INV_39\, \AFLSDF_INV_40\, 
        \AFLSDF_INV_41\, \AFLSDF_INV_42\, \AFLSDF_INV_43\, 
        \AFLSDF_INV_44\, \AFLSDF_INV_45\, \AFLSDF_INV_46\, 
        \AFLSDF_INV_47\, \AFLSDF_INV_48\, \AFLSDF_INV_49\, 
        \AFLSDF_INV_50\, \AFLSDF_INV_51\, \AFLSDF_INV_52\, 
        \AFLSDF_INV_53\, \AFLSDF_INV_54\, \AFLSDF_INV_55\, 
        \AFLSDF_INV_56\, \AFLSDF_INV_57\, \AFLSDF_INV_58\, 
        \AFLSDF_INV_59\, \AFLSDF_INV_60\, \AFLSDF_INV_61\, 
        \AFLSDF_INV_62\, \AFLSDF_INV_63\, \AFLSDF_INV_64\, 
        \AFLSDF_INV_65\, \AFLSDF_INV_66\, \AFLSDF_INV_67\, 
        \AFLSDF_INV_68\, \AFLSDF_INV_69\, \AFLSDF_INV_70\, 
        \AFLSDF_INV_71\, \AFLSDF_INV_72\, \AFLSDF_INV_73\, 
        \AFLSDF_INV_74\, \AFLSDF_INV_75\, \AFLSDF_INV_76\, 
        \AFLSDF_INV_77\, \AFLSDF_INV_78\, \AFLSDF_INV_79\, 
        \AFLSDF_INV_80\, \AFLSDF_INV_81\, \AFLSDF_INV_82\, 
        \AFLSDF_INV_83\, \AFLSDF_INV_84\, \AFLSDF_INV_85\, 
        \AFLSDF_INV_86\, \AFLSDF_INV_87\, \AFLSDF_INV_88\, 
        \AFLSDF_INV_89\, \AFLSDF_INV_90\, \AFLSDF_INV_91\, 
        \AFLSDF_INV_92\, \AFLSDF_INV_93\, \AFLSDF_INV_94\, 
        \AFLSDF_INV_95\, \AFLSDF_INV_96\, \AFLSDF_INV_97\, 
        \AFLSDF_INV_98\, \AFLSDF_INV_99\, \AFLSDF_INV_100\, 
        \AFLSDF_INV_101\, \AFLSDF_INV_102\, \AFLSDF_INV_103\, 
        \AFLSDF_INV_104\, \AFLSDF_INV_105\, \AFLSDF_INV_106\, 
        \AFLSDF_INV_107\, \AFLSDF_INV_108\, \AFLSDF_INV_109\, 
        \AFLSDF_INV_110\, \AFLSDF_INV_111\, \AFLSDF_INV_112\
         : std_logic;
    signal GND_power_net1 : std_logic;
    signal VCC_power_net1 : std_logic;
    signal nc228, nc203, nc265, nc216, nc194, nc151, nc23, nc440, 
        nc175, nc393, nc250, nc411, nc58, nc379, nc116, nc74, 
        nc133, nc420, nc238, nc167, nc84, nc39, nc72, nc256, 
        nc212, nc205, nc82, nc367, nc145, nc181, nc160, nc57, 
        nc430, nc349, nc156, nc395, nc280, nc125, nc211, nc73, 
        nc107, nc408, nc329, nc66, nc83, nc9, nc252, nc171, nc54, 
        nc286, nc307, nc135, nc41, nc100, nc404, nc270, nc339, 
        nc52, nc251, nc186, nc29, nc269, nc118, nc412, nc60, 
        nc141, nc311, nc276, nc193, nc214, nc298, nc282, nc240, 
        nc45, nc53, nc121, nc176, nc419, nc360, nc220, nc158, 
        nc281, nc209, nc427, nc246, nc368, nc351, nc162, nc11, 
        nc272, nc131, nc364, nc254, nc267, nc96, nc79, nc441, 
        nc226, nc146, nc230, nc89, nc119, nc48, nc437, nc271, 
        nc213, nc421, nc366, nc300, nc126, nc195, nc188, nc242, 
        nc15, nc399, nc308, nc236, nc102, nc381, nc304, nc3, 
        nc207, nc47, nc90, nc284, nc222, nc159, nc431, nc136, 
        nc241, nc253, nc178, nc306, nc215, nc59, nc362, nc221, 
        nc371, nc232, nc274, nc18, nc44, nc117, nc418, nc189, 
        nc164, nc148, nc42, nc231, nc191, nc255, nc442, nc283, 
        nc363, nc341, nc317, nc290, nc17, nc2, nc406, nc302, 
        nc110, nc128, nc414, nc244, nc422, nc321, nc43, nc179, 
        nc157, nc36, nc224, nc296, nc273, nc61, nc104, nc138, 
        nc14, nc432, nc357, nc285, nc429, nc405, nc303, nc150, 
        nc365, nc331, nc196, nc234, nc149, nc12, nc219, nc30, 
        nc243, nc187, nc65, nc7, nc292, nc439, nc129, nc275, nc8, 
        nc223, nc13, nc387, nc305, nc180, nc26, nc291, nc177, 
        nc139, nc310, nc259, nc403, nc245, nc233, nc163, nc318, 
        nc268, nc112, nc68, nc49, nc377, nc314, nc217, nc170, 
        nc91, nc225, nc5, nc20, nc198, nc147, nc350, nc316, nc391, 
        nc67, nc289, nc358, nc294, nc152, nc127, nc103, nc428, 
        nc235, nc76, nc347, nc208, nc354, nc140, nc257, nc86, 
        nc95, nc327, nc120, nc424, nc165, nc356, nc279, nc137, 
        nc438, nc64, nc400, nc19, nc380, nc369, nc416, nc312, 
        nc70, nc388, nc182, nc62, nc337, nc199, nc80, nc130, 
        nc434, nc384, nc287, nc98, nc293, nc249, nc114, nc56, 
        nc370, nc105, nc386, nc63, nc415, nc352, nc313, nc309, 
        nc378, nc172, nc229, nc374, nc277, nc97, nc161, nc31, 
        nc340, nc295, nc154, nc376, nc50, nc260, nc239, nc353, 
        nc348, nc142, nc320, nc344, nc315, nc382, nc247, nc94, 
        nc197, nc328, nc122, nc266, nc35, nc324, nc4, nc227, nc92, 
        nc101, nc413, nc346, nc330, nc397, nc184, nc200, nc190, 
        nc166, nc372, nc407, nc355, nc338, nc326, nc132, nc383, 
        nc334, nc21, nc237, nc93, nc262, nc69, nc206, nc174, nc38, 
        nc113, nc336, nc218, nc401, nc342, nc373, nc106, nc261, 
        nc25, nc1, nc385, nc426, nc322, nc299, nc37, nc410, nc202, 
        nc144, nc153, nc46, nc258, nc343, nc71, nc124, nc436, 
        nc332, nc81, nc375, nc201, nc168, nc425, nc323, nc390, 
        nc34, nc28, nc361, nc115, nc264, nc398, nc192, nc319, 
        nc134, nc394, nc32, nc40, nc297, nc99, nc75, nc183, nc435, 
        nc345, nc333, nc288, nc85, nc27, nc108, nc396, nc402, 
        nc325, nc16, nc155, nc51, nc301, nc33, nc443, nc359, 
        nc204, nc173, nc278, nc169, nc423, nc78, nc263, nc335, 
        nc24, nc409, nc88, nc111, nc55, nc10, nc22, nc392, nc210, 
        nc185, nc143, nc433, nc417, nc248, nc389, nc77, nc6, 
        nc109, nc87, nc123 : std_logic;

    for all : sdf_IOPAD_TRI
	Use entity work.sdf_IOPAD_TRI(DEF_ARCH);
    for all : sdf_IOPAD_IN
	Use entity work.sdf_IOPAD_IN(DEF_ARCH);
begin 

    ADLIB_GND0 <= GND_power_net1;
    AFLSDF_GND <= GND_power_net1;
    ADLIB_VCC1 <= VCC_power_net1;
    AFLSDF_VCC <= VCC_power_net1;

    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_229\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_193\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_41_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_0\, ADn => ADLIB_GND0, SLn
         => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_41_set_Z\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_36\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[30]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_36_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[4]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[4]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[4]\, D => 
        \MemorySynchronizer_0/un5_resettimercounter_m[28]\, Y => 
        \MemorySynchronizer_0/resettimercounter_9[4]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_10\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[10]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[10]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_9\, S => 
        \MemorySynchronizer_0/temp_1[10]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_10\, CC => 
        NET_CC_CONFIG229, P => NET_CC_CONFIG227, UB => 
        NET_CC_CONFIG228);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1[20]\ : 
        CFG4
      generic map(INIT => x"F3FB")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => \MemorySynchronizer_0/un151_in_enable\, C => 
        \MemorySynchronizer_0/N_2328\, D => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, Y
         => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[14]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[14]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[18]\, Y
         => \MemorySynchronizer_0/N_1077\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_14\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[14]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_13_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_14_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_14_Z\, CC
         => NET_CC_CONFIG767, P => NET_CC_CONFIG765, UB => 
        NET_CC_CONFIG766);
    
    \MemorySynchronizer_0/TimeStampGen/counter[20]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[20]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[20]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_12\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[12]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_11_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_12_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_12_Z\, CC
         => NET_CC_CONFIG761, P => NET_CC_CONFIG759, UB => 
        NET_CC_CONFIG760);
    
    \MemorySynchronizer_0/un104_in_enable_cry_3\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[3]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[3]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_2_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_3_Z\, CC => 
        NET_CC_CONFIG832, P => NET_CC_CONFIG830, UB => 
        NET_CC_CONFIG831);
    
    \STAMP_0/async_prescaler_count_5[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/un1_async_prescaler_count\, B => 
        \STAMP_0/un5_async_prescaler_count_cry_6_S\, Y => 
        \STAMP_0/async_prescaler_count_5_Z[6]\);
    
    \STAMP_0/dummy[18]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_1\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[18]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_25\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[18]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[18]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[14]\, Y
         => \MemorySynchronizer_0/N_1073\);
    
    \STAMP_0/status_async_cycles_lm_0[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/status_async_cycles_3_sqmuxa\, B => 
        \STAMP_0/status_async_cycles_s[1]\, C => 
        \STAMP_0/status_async_cycles_1_sqmuxa_Z\, Y => 
        \STAMP_0/status_async_cycles_lm[1]\);
    
    \STAMP_0/spi/tx_buffer[14]\ : SLE
      port map(D => \STAMP_0/spi/N_121\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[14]\);
    
    \MemorySynchronizer_0/un1_nreset_34_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_53_i_i_a2_Z\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_34_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_34_rs_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_6[28]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[28]\, 
        B => \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2567\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1168\);
    
    AFLSDF_INV_36 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_36\);
    
    \STAMP_0/spi/tx_buffer[6]\ : SLE
      port map(D => \STAMP_0/spi/N_130\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[6]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[6]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[6]\, B => 
        \sb_sb_0_STAMP_PWDATA[6]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[6]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_19\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[19]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_18_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[13]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_19_Z\, CC
         => NET_CC_CONFIG354, P => NET_CC_CONFIG352, UB => 
        NET_CC_CONFIG353);
    
    \STAMP_0/spi/count_cry[29]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[29]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[28]\, S => 
        \STAMP_0/spi/count_s[29]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[29]\, CC => NET_CC_CONFIG1012, P
         => NET_CC_CONFIG1010, UB => NET_CC_CONFIG1011);
    
    \MemorySynchronizer_0/un1_nreset_6_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_36_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_6_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_6_rs_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4[16]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \MemorySynchronizer_0/un104_in_enable_16\, B
         => \MemorySynchronizer_0/SynchStatusReg2_Z[16]\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2594\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[16]\);
    
    \STAMP_0/PRDATA[28]\ : SLE
      port map(D => \STAMP_0/N_678\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_2\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[28]\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => OPEN, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[12]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[12]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[11]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[12]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[12]\, CC
         => NET_CC_CONFIG42, P => NET_CC_CONFIG40, UB => 
        NET_CC_CONFIG41);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_41_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_3\, ADn => ADLIB_GND0, SLn
         => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_41_set_Z\);
    
    \STAMP_0/un1_async_state_0_sqmuxa\ : CFG4
      generic map(INIT => x"FFBA")

      port map(A => \STAMP_0/request_resync_0_sqmuxa\, B => 
        sb_sb_0_STAMP_PENABLE, C => 
        \STAMP_0/async_state_0_sqmuxa_1_1_Z\, D => 
        \STAMP_0/async_state_0_sqmuxa_Z\, Y => 
        \STAMP_0/un1_async_state_0_sqmuxa_i\);
    
    \STAMP_0/dummy[26]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_4\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[26]\);
    
    \STAMP_0/PRDATA[9]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[9]\);
    
    \STAMP_0/delay_counter_cry[24]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[24]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[23]\, S
         => \STAMP_0/delay_counter_s[24]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[24]\, CC => NET_CC_CONFIG467, 
        P => NET_CC_CONFIG465, UB => NET_CC_CONFIG466);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB7\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\);
    
    \MemorySynchronizer_0/waitingtimercounter[8]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_58_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[8]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_56\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17]\, 
        IPC => OPEN);
    
    AFLSDF_INV_51 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_31\, Y => 
        \AFLSDF_INV_51\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_15\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[15]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_14_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_15_Z\, CC => 
        NET_CC_CONFIG868, P => NET_CC_CONFIG866, UB => 
        NET_CC_CONFIG867);
    
    AFLSDF_INV_90 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_49_Z\, Y => 
        \AFLSDF_INV_90\);
    
    \ENABLE_MEMORY_LED_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => ENABLE_MEMORY_LED, D => 
        \ENABLE_MEMORY_LED_obuf/U0/DOUT\, E => 
        \ENABLE_MEMORY_LED_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_43\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[17]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_43_Z\);
    
    \MemorySynchronizer_0/MemorySyncState_RNIFKGB[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ENABLE_MEMORY_LED_c, B => 
        \MemorySynchronizer_0/MemorySyncState_Z[3]\, Y => 
        \MemorySynchronizer_0/N_140_1_i\);
    
    \STAMP_0/status_async_cycles[2]\ : SLE
      port map(D => \STAMP_0/status_async_cycles_lm[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/status_async_cycles_1_sqmuxa_1_i_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[5]\);
    
    \STAMP_0/un1_presetn_inv_2_i_0\ : CFG4
      generic map(INIT => x"C444")

      port map(A => \STAMP_0/N_219\, B => debug_led_net_0, C => 
        \STAMP_0/config_Z[30]\, D => \STAMP_0/N_333\, Y => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_277\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4]\, 
        IPC => OPEN);
    
    \STAMP_0/async_prescaler_count[4]\ : SLE
      port map(D => \STAMP_0/un5_async_prescaler_count_cry_4_S\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[4]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_76\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17]\, 
        IPC => OPEN);
    
    \STAMP_0/measurement_dms2[9]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[41]\);
    
    \MemorySynchronizer_0/resettimercounter[23]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_10_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[23]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_99\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[6]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un5_resettimercounter_s_31\ : ARI1_CC
      generic map(INIT => x"45500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[31]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_30_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_s_31_S\, 
        Y => OPEN, FCO => OPEN, CC => NET_CC_CONFIG818, P => 
        NET_CC_CONFIG816, UB => NET_CC_CONFIG817);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_21\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[23]\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[21]\, C => 
        \MemorySynchronizer_0/waitingtimercounter_Z[20]\, D => 
        \MemorySynchronizer_0/waitingtimercounter_Z[13]\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_21_Z\);
    
    \STAMP_0/spi/count_s_389_CC_0\ : CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => CI_TO_CO920, P(0) => 
        ADLIB_VCC1, P(1) => ADLIB_VCC1, P(2) => ADLIB_VCC1, P(3)
         => ADLIB_VCC1, P(4) => ADLIB_VCC1, P(5) => ADLIB_VCC1, 
        P(6) => ADLIB_VCC1, P(7) => ADLIB_VCC1, P(8) => 
        ADLIB_VCC1, P(9) => ADLIB_VCC1, P(10) => ADLIB_GND0, 
        P(11) => NET_CC_CONFIG923, UB(0) => ADLIB_VCC1, UB(1) => 
        ADLIB_VCC1, UB(2) => ADLIB_VCC1, UB(3) => ADLIB_VCC1, 
        UB(4) => ADLIB_VCC1, UB(5) => ADLIB_VCC1, UB(6) => 
        ADLIB_VCC1, UB(7) => ADLIB_VCC1, UB(8) => ADLIB_VCC1, 
        UB(9) => ADLIB_VCC1, UB(10) => ADLIB_GND0, UB(11) => 
        NET_CC_CONFIG924, CC(0) => nc228, CC(1) => nc203, CC(2)
         => nc265, CC(3) => nc216, CC(4) => nc194, CC(5) => nc151, 
        CC(6) => nc23, CC(7) => nc440, CC(8) => nc175, CC(9) => 
        nc393, CC(10) => nc250, CC(11) => NET_CC_CONFIG925);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[4]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[4]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[27]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB0_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[27]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[2]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[2]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[2]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[2]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[2]\);
    
    \STAMP_0/status_dms2_newVal\ : SLE
      port map(D => \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_1\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, 
        EN => \STAMP_0/un1_new_avail_0_sqmuxa_3_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[14]\);
    
    \MemorySynchronizer_0/un1_nreset_54_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[12]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_54_i\);
    
    \STAMP_0/spi/rx_buffer[7]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[7]\);
    
    \STAMP_0/measurement_dms2[10]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[42]\);
    
    \STAMP_0/delay_counter_cry[15]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[15]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[14]\, S
         => \STAMP_0/delay_counter_s[15]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[15]\, CC => NET_CC_CONFIG440, 
        P => NET_CC_CONFIG438, UB => NET_CC_CONFIG439);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[2]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[2]\, B => 
        \sb_sb_0_STAMP_PWDATA[2]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[2]\);
    
    \STAMP_0/config[30]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[30]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[30]\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_s_387\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[0]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => ADLIB_VCC1, S => OPEN, Y => OPEN, 
        FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_s_387_FCO\, CC
         => NET_CC_CONFIG6, P => NET_CC_CONFIG4, UB => 
        NET_CC_CONFIG5);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB12\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => OPEN, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB12_rgbr_net_1\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_42\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net\, IPC
         => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_259\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19]\, 
        IPC => OPEN);
    
    \STAMP_0/dummy[21]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_5\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[21]\);
    
    \MemorySynchronizer_0/MemorySyncState[3]\ : SLE
      port map(D => \MemorySynchronizer_0/MemorySyncState_ns[2]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, 
        EN => ENABLE_MEMORY_LED_c, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/MemorySyncState_Z[3]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[6]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[6]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1[26]\, Y => 
        \MemorySynchronizer_0/N_1085\);
    
    \STAMP_0/spi/count[1]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[1]\);
    
    \STAMP_0/spi_tx_data[10]\ : SLE
      port map(D => \STAMP_0/un1_pwdata_Z[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[10]\);
    
    \STAMP_0/delay_counter_lm_0[20]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[20]\, Y => 
        \STAMP_0/delay_counter_lm[20]\);
    
    \STAMP_0/spi/count_lm_0[1]\ : CFG4
      generic map(INIT => x"D8CC")

      port map(A => \STAMP_0/spi/un7_count_NE_i\, B => 
        \STAMP_0/spi/count_0_sqmuxa\, C => 
        \STAMP_0/spi/count_s[1]\, D => \STAMP_0/spi/state_Z[0]\, 
        Y => \STAMP_0/spi/count_lm[1]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_30\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/N_2536_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_6\, ADn => ADLIB_GND0, SLn
         => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_2536_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_178\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[7]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => \MemorySynchronizer_0/N_1182\, B => 
        \MemorySynchronizer_0/N_2575\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[7]\, D => 
        \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[7]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_41_set_RNIPMAM\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_41_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[4]\, C
         => \MemorySynchronizer_0/un1_nreset_4_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[4]\);
    
    \STAMP_0/spi/count_lm_0[16]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[16]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[16]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[0]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB0_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[0]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_261\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_47_i_i_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[26]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_47_i_i_a2_Z\);
    
    \MemorySynchronizer_0/resynctimercounter[26]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1096\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[26]\);
    
    \MemorySynchronizer_0/resettimercounter_RNI22C41[16]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_44_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[16]\, C => 
        \MemorySynchronizer_0/un1_nreset_17_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[16]\);
    
    AFLSDF_INV_62 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_62\);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_19\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[28]\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[26]\, C => 
        \MemorySynchronizer_0/waitingtimercounter_Z[18]\, D => 
        \MemorySynchronizer_0/waitingtimercounter_Z[16]\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_19_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_24[10]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[3]\, D => \sb_sb_0_STAMP_PADDR[4]\, 
        Y => \MemorySynchronizer_0/N_2580\);
    
    \STAMP_0/spi/count[20]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[20]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[21]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_21\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[21]\, 
        C => \MemorySynchronizer_0/N_1497\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[21]\);
    
    \MemorySynchronizer_0/un1_nreset_42_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[24]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_42_i\);
    
    \STAMP_0/spi/tx_buffer_RNO[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[3]\, B => 
        \STAMP_0/spi/tx_buffer_Z[2]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_136\);
    
    \STAMP_0/delay_counter_lm_0[21]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[21]\, Y => 
        \STAMP_0/delay_counter_lm[21]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_283\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10]\, 
        IPC => OPEN);
    
    \STAMP_0/delay_counter[18]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[18]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[4]\ : SLE
      port map(D => \MemorySynchronizer_0/temp_1[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[4]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_25[20]\ : 
        CFG4
      generic map(INIT => x"1000")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[10]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[28]\, C => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_19_Z[20]\, 
        D => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_10_Z[20]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_25_Z[20]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_1\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[1]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[1]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_0_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_1_Z\, CC => 
        NET_CC_CONFIG826, P => NET_CC_CONFIG824, UB => 
        NET_CC_CONFIG825);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[19]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[19]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[13]\, Y
         => \MemorySynchronizer_0/N_1072\);
    
    \STAMP_0/spi/count_cry[10]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[10]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[9]\, S => 
        \STAMP_0/spi/count_s[10]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[10]\, CC => NET_CC_CONFIG955, P
         => NET_CC_CONFIG953, UB => NET_CC_CONFIG954);
    
    \STAMP_0/delay_counter_RNIUVPA[24]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \STAMP_0/delay_counter_Z[27]\, B => 
        \STAMP_0/delay_counter_Z[26]\, C => 
        \STAMP_0/delay_counter_Z[25]\, D => 
        \STAMP_0/delay_counter_Z[24]\, Y => 
        \STAMP_0/N_517_i_0_a2_20\);
    
    \MemorySynchronizer_0/SynchStatusReg2[21]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[21]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_199\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[12]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_72\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[12]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[12]\, 
        D => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[12]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_55_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_7\, ADn => ADLIB_GND0, SLn
         => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_55_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_247\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7]\, IPC
         => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_195\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_56\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[6]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_ResetTimerValueReg_56_Z\);
    
    \MemorySynchronizer_0/numberofnewavails[0]\ : SLE
      port map(D => \MemorySynchronizer_0/ConfigReg_Z[0]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/numberofnewavails_0_sqmuxa\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/numberofnewavails_Z[0]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_11\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[11]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_10_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[11]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_11_Z\, 
        CC => NET_CC_CONFIG137, P => NET_CC_CONFIG135, UB => 
        NET_CC_CONFIG136);
    
    \MemorySynchronizer_0/PRDATA[27]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[27]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[27]\);
    
    \STAMP_0/spi/count[24]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[24]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_15[19]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_18_0_Z[19]\, B
         => \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[5]\, Y => 
        \MemorySynchronizer_0/N_2572\);
    
    \STAMP_0/delay_counter[22]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[22]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[14]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[14]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[14]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_53_i_i_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[0]\, B => NN_1, 
        Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_53_i_i_a2_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[6]\ : CFG4
      generic map(INIT => x"CCA0")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_m_0_0[6]\, B => 
        \sb_sb_0_STAMP_PWDATA[6]\, C => ENABLE_MEMORY_LED_c, D
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[6]\);
    
    \STAMP_0/un1_spi_rx_data_2[13]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_596\, B => \STAMP_0/N_630\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_663\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_14\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[14]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_13_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_14_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_14_Z\, 
        CC => NET_CC_CONFIG669, P => NET_CC_CONFIG667, UB => 
        NET_CC_CONFIG668);
    
    \STAMP_0/spi/count[7]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[7]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_45\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_182\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_62_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_32\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_62_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_62_rs_Z\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[23]\ : SLE
      port map(D => \STAMP_0_data_frame[55]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[23]\);
    
    \STAMP_0/spi/rx_buffer[9]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[9]\);
    
    \MemorySynchronizer_0/un1_nreset_48\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[7]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_48_i\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[5]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[5]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[5]\, C => 
        \MemorySynchronizer_0/un104_in_enable_5\, D => 
        \MemorySynchronizer_0/N_1204_1\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[5]\);
    
    \MemorySynchronizer_0/PRDATA[14]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[14]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[14]\);
    
    \STAMP_0/PRDATA[24]\ : SLE
      port map(D => \STAMP_0/N_674\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_8\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[24]\);
    
    \MemorySynchronizer_0/un1_nreset_22_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[22]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_22_i\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbl_net_1\, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\);
    
    \STAMP_0/spi_tx_data[8]\ : SLE
      port map(D => \STAMP_0/N_290_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[8]\);
    
    \STAMP_0/spi_request_for[0]\ : SLE
      port map(D => \STAMP_0/N_567_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_4_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_request_for_Z[0]\);
    
    AFLSDF_INV_9 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_9\);
    
    \STAMP_0/un5_async_prescaler_count_s_1_391_CC_1\ : CC_CONFIG
      port map(CI => CI_TO_CO477, CO => OPEN, P(0) => 
        NET_CC_CONFIG487, P(1) => NET_CC_CONFIG490, P(2) => 
        NET_CC_CONFIG493, P(3) => NET_CC_CONFIG496, P(4) => 
        NET_CC_CONFIG499, P(5) => NET_CC_CONFIG502, P(6) => 
        NET_CC_CONFIG505, P(7) => NET_CC_CONFIG508, P(8) => 
        NET_CC_CONFIG511, P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, 
        P(11) => ADLIB_VCC1, UB(0) => NET_CC_CONFIG488, UB(1) => 
        NET_CC_CONFIG491, UB(2) => NET_CC_CONFIG494, UB(3) => 
        NET_CC_CONFIG497, UB(4) => NET_CC_CONFIG500, UB(5) => 
        NET_CC_CONFIG503, UB(6) => NET_CC_CONFIG506, UB(7) => 
        NET_CC_CONFIG509, UB(8) => NET_CC_CONFIG512, UB(9) => 
        ADLIB_VCC1, UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, 
        CC(0) => NET_CC_CONFIG489, CC(1) => NET_CC_CONFIG492, 
        CC(2) => NET_CC_CONFIG495, CC(3) => NET_CC_CONFIG498, 
        CC(4) => NET_CC_CONFIG501, CC(5) => NET_CC_CONFIG504, 
        CC(6) => NET_CC_CONFIG507, CC(7) => NET_CC_CONFIG510, 
        CC(8) => NET_CC_CONFIG513, CC(9) => nc411, CC(10) => nc58, 
        CC(11) => nc379);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[21]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_88\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[21]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[21]\, 
        D => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[21]\);
    
    \STAMP_0/un1_spi_rx_data_1[5]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[37]\, B => 
        \STAMP_0/dummy_Z[5]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_622\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_285\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_148\ : 
        IP_INTERFACE
      port map(A => RXSM_SOE_c, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/ConfigReg[10]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[10]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_4\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[4]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[4]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_3_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_4_Z\, CC => 
        NET_CC_CONFIG835, P => NET_CC_CONFIG833, UB => 
        NET_CC_CONFIG834);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_278\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5]\, 
        IPC => OPEN);
    
    \STAMP_0/delay_counter[20]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[20]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_18\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[18]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_17_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[14]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_18_Z\, CC
         => NET_CC_CONFIG351, P => NET_CC_CONFIG349, UB => 
        NET_CC_CONFIG350);
    
    \STAMP_0/measurement_dms2[4]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[36]\);
    
    \MemorySynchronizer_0/SynchStatusReg_152_sn.m3_1_0_o2\ : CFG4
      generic map(INIT => x"3337")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => ENABLE_MEMORY_LED_c, C => 
        \MemorySynchronizer_0/MemorySyncState_Z[0]\, D => 
        \MemorySynchronizer_0/MemorySyncState_Z[2]\, Y => 
        \MemorySynchronizer_0/un1_enabletimestampgen2_2_sn\);
    
    \MemorySynchronizer_0/ReadInterrupt_0_sqmuxa_2_i_0_a2_1\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/N_2567\, B => 
        \MemorySynchronizer_0/N_2586\, C => 
        \MemorySynchronizer_0/APBState_Z[1]\, D => 
        \sb_sb_0_STAMP_PWDATA[29]\, Y => 
        \MemorySynchronizer_0/N_191\);
    
    \MemorySynchronizer_0/PRDATA[0]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[0]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[0]\);
    
    \STAMP_0/un1_spi_rx_data_1[16]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[48]\, B => 
        \STAMP_0/dummy_Z[16]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_633\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[20]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[20]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[20]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[12]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[20]\);
    
    \STAMP_0/PRDATA[0]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[0]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_8\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_9\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_7_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[9]\, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_8_Z\, 
        CC => NET_CC_CONFIG1047, P => NET_CC_CONFIG1045, UB => 
        NET_CC_CONFIG1046);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_69\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_o2[30]\ : 
        CFG3
      generic map(INIT => x"FE")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => \MemorySynchronizer_0/MemorySyncState_Z[5]\, C => 
        \MemorySynchronizer_0/MemorySyncState_Z[2]\, Y => 
        \MemorySynchronizer_0/N_2315\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_1\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net\, IPB
         => OPEN, IPC => OPEN);
    
    \STAMP_0/config[0]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[0]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_196\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12]\, 
        IPC => OPEN);
    
    \AND2_0_RNIKOS1/U0_RGB1_RGB1\ : RGB_NG
      port map(An => \AND2_0_RNIKOS1/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[25]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[25]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[27]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[25]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[15]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[15]\, B => 
        \sb_sb_0_Memory_PRDATA[15]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[30]\ : SLE
      port map(D => \STAMP_0_data_frame[30]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[30]\);
    
    \STAMP_0/spi/count_lm_0[19]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[19]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[19]\);
    
    \STAMP_0/dummy[17]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_9\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[17]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[16]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_16\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_9\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[9]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_8_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[9]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_9_Z\, 
        CC => NET_CC_CONFIG131, P => NET_CC_CONFIG129, UB => 
        NET_CC_CONFIG130);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_16\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[16]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_15_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_16_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_16_Z\, CC
         => NET_CC_CONFIG773, P => NET_CC_CONFIG771, UB => 
        NET_CC_CONFIG772);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_19_Z\, B
         => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_18_Z\, 
        C => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_31_Z\, 
        D => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_27_Z\, 
        Y => \MemorySynchronizer_0/un41_in_enable_i_0\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_30\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[30]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[30]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_29\, S => 
        \MemorySynchronizer_0/temp_1[30]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_30_FCNET1\, 
        CC => NET_CC_CONFIG289, P => NET_CC_CONFIG287, UB => 
        NET_CC_CONFIG288);
    
    \MemorySynchronizer_0/un1_nreset_15_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_42_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_15_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_15_rs_Z\);
    
    \MemorySynchronizer_0/un1_nreset_2_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[3]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_2_i\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[9]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_9_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[23]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[21]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_21\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[21]\ : SLE
      port map(D => \STAMP_0_data_frame[53]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[21]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_123\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_18\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[18]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_17_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[18]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_18_Z\, 
        CC => NET_CC_CONFIG158, P => NET_CC_CONFIG156, UB => 
        NET_CC_CONFIG157);
    
    \MemorySynchronizer_0/waitingtimercounter_RNI1B6R[17]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_61_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[17]\, C
         => \MemorySynchronizer_0/un1_nreset_24_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[17]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_38_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_10\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_38_set_Z\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_11\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[11]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_10_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_11_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_11_Z\, 
        CC => NET_CC_CONFIG660, P => NET_CC_CONFIG658, UB => 
        NET_CC_CONFIG659);
    
    \MemorySynchronizer_0/N_1978_i_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_11\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_1978_i_set_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[6]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_6_S\, 
        Y => \MemorySynchronizer_0/N_1541\);
    
    \MemorySynchronizer_0/TimeStampReg[7]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[7]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[7]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[7]\ : SLE
      port map(D => \STAMP_0_data_frame[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[7]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[22]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[22]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1069\, Y => 
        \MemorySynchronizer_0/N_1100\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[16]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_16_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[16]\);
    
    \STAMP_0/spi/mosi_1_1_0_0_a2_2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \STAMP_0/spi/assert_data_Z\, B => 
        \STAMP_0/spi/clk_toggles_Z[5]\, C => 
        \STAMP_0/spi/state_Z[0]\, D => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/mosi_1_1_2\);
    
    \STAMP_0/spi/un7_count_NE_16\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \STAMP_0/spi/count_Z[19]\, B => 
        \STAMP_0/spi/count_Z[18]\, C => \STAMP_0/spi/count_Z[17]\, 
        D => \STAMP_0/spi/count_Z[16]\, Y => 
        \STAMP_0/spi/un7_count_NE_16_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[20]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[20]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[20]\, D
         => \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[20]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[14]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[14]\);
    
    \MemorySynchronizer_0/resettimercounter[14]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_7_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[14]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[2]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[2]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[2]\, D => 
        \MemorySynchronizer_0/un5_resettimercounter_m[30]\, Y => 
        \MemorySynchronizer_0/resettimercounter_9[2]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_o2_1[4]\ : 
        CFG4
      generic map(INIT => x"4505")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[5]\, 
        B => STAMP_0_new_avail, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, Y
         => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_o2_1_0[4]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_33_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[16]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_33\);
    
    \STAMP_0/apb_is_atomic\ : SLE
      port map(D => \sb_sb_0_STAMP_PADDR[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/apb_is_atomic_0_sqmuxa\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/apb_is_atomic_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_15[28]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \MemorySynchronizer_0/N_2576\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, Y => 
        \MemorySynchronizer_0/N_2597\);
    
    \STAMP_0/spi/tx_buffer_RNO[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[9]\, B => 
        \STAMP_0/spi/tx_buffer_Z[8]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_126\);
    
    \STAMP_0/async_prescaler_count_5[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/un1_async_prescaler_count\, B => 
        \STAMP_0/un5_async_prescaler_count_cry_2_S\, Y => 
        \STAMP_0/async_prescaler_count_5_Z[2]\);
    
    \MemorySynchronizer_0/ReadInterrupt_RNO\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \MemorySynchronizer_0/N_2567\, B => 
        \MemorySynchronizer_0/N_2586\, C => 
        \MemorySynchronizer_0/APBState_Z[1]\, D => 
        \sb_sb_0_STAMP_PWDATA[29]\, Y => 
        \MemorySynchronizer_0/N_191_i\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_21\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/N_1090\, B => 
        \MemorySynchronizer_0/N_1074\, C => 
        \MemorySynchronizer_0/N_1073\, D => 
        \MemorySynchronizer_0/N_1072\, Y => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_21_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[25]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[25]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[25]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[9]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[9]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[22]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[22]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_29\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[29]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[29]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_28\, S => 
        \MemorySynchronizer_0/temp_1[29]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_29\, CC => 
        NET_CC_CONFIG286, P => NET_CC_CONFIG284, UB => 
        NET_CC_CONFIG285);
    
    \STAMP_0/dummy[14]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_12\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[14]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_40\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[20]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_40_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[25]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_25_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[7]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[23]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[23]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[23]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[23]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[23]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[23]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_46_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_13\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_46_set_Z\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_45\ : ARI1_CC
      generic map(INIT => x"62100")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_30\, C => 
        \MemorySynchronizer_0/un104_in_enable_axb_31\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[30]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[14]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_I_45_FCNET1\, CC
         => NET_CC_CONFIG583, P => NET_CC_CONFIG581, UB => 
        NET_CC_CONFIG582);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_2\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_3\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_1_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[3]\, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_2_Z\, 
        CC => NET_CC_CONFIG1029, P => NET_CC_CONFIG1027, UB => 
        NET_CC_CONFIG1028);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[25]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[25]\, B => 
        \MemorySynchronizer_0/un104_in_enable_25\, C => 
        \MemorySynchronizer_0/N_2574\, D => 
        \MemorySynchronizer_0/N_2577\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[25]\);
    
    \STAMP_0/component_state[3]\ : SLE
      port map(D => \STAMP_0/component_state_ns[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/component_state_Z[3]\);
    
    \MemorySynchronizer_0/un1_nreset_56_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_56_i_i_a2_Z\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_56_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_56_rs_Z\);
    
    \sb_sb_0/CCC_0/GL1_INST\ : GB_NG
      port map(An => \AFLSDF_INV_14\, ENn => ADLIB_GND0, YNn => 
        OPEN, YSn => \sb_sb_0/CCC_0/GL1_INST/U0_YNn_GSouth\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_11\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_12\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_10_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[12]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_11_Z\, CC
         => NET_CC_CONFIG1056, P => NET_CC_CONFIG1054, UB => 
        NET_CC_CONFIG1055);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_2\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0]\, B
         => ADLIB_VCC1, C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0]\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/un52_paddr_2_0_a2\ : CFG2
      generic map(INIT => x"1")

      port map(A => \sb_sb_0_STAMP_PADDR[8]\, B => 
        \sb_sb_0_STAMP_PADDR[4]\, Y => \STAMP_0/un52_paddr_2_Z\);
    
    \STAMP_0/un1_component_state_9_i_o2_1\ : CFG4
      generic map(INIT => x"F8FF")

      port map(A => \STAMP_0/N_109_i\, B => \STAMP_0/N_238\, C
         => \STAMP_0/config_Z[31]\, D => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_215\);
    
    \MemorySynchronizer_0/waitingtimercounter_RNIOJ601[22]\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_40_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[22]\, C
         => \MemorySynchronizer_0/un1_nreset_22_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[22]\);
    
    \STAMP_0/spi/rx_data[2]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB0_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[2]\);
    
    \STAMP_0/delay_counter_lm_0[15]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[15]\, Y => 
        \STAMP_0/delay_counter_lm[15]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_248\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, B
         => \MemorySynchronizer_0/resettimercounter_Z[6]\, Y => 
        \MemorySynchronizer_0/resettimercounter_m[6]\);
    
    \MemorySynchronizer_0/ConfigReg[29]\ : SLE
      port map(D => \MemorySynchronizer_0/N_2305_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/un1_APBState_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[29]\);
    
    \STAMP_0/config[2]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[2]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_15\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[15]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_14_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_15_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_15_Z\, CC
         => NET_CC_CONFIG770, P => NET_CC_CONFIG768, UB => 
        NET_CC_CONFIG769);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[13]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[13]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[13]\, C => 
        \MemorySynchronizer_0/N_2596\, D => 
        \MemorySynchronizer_0/N_2595\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[13]\);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB4\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[8]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[8]\, B => 
        \MemorySynchronizer_0/N_2567\, C => 
        \MemorySynchronizer_0/N_2586\, Y => 
        \MemorySynchronizer_0/N_1245\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_92\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_ERRF_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_50\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[5]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_50_i\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_10\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[10]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_9_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_10_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_10_Z\, 
        CC => NET_CC_CONFIG657, P => NET_CC_CONFIG655, UB => 
        NET_CC_CONFIG656);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[14]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[14]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[14]\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[14]\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[14]\);
    
    \STAMP_0/un1_spi_rx_data_2[10]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_593\, B => \STAMP_0/N_627\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_660\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_0\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[0]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => ADLIB_GND0, S => OPEN, Y => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_Y\, 
        FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_Z\, 
        CC => NET_CC_CONFIG104, P => NET_CC_CONFIG102, UB => 
        NET_CC_CONFIG103);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_18\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[23]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[30]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30]\, 
        IPC => OPEN);
    
    \STAMP_0/delay_counter[25]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[25]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_2\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[2]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_1_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[30]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_2_Z\, CC
         => NET_CC_CONFIG303, P => NET_CC_CONFIG301, UB => 
        NET_CC_CONFIG302);
    
    \MemorySynchronizer_0/un1_nreset_35_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_42\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_35_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_35_rs_Z\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[5]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[5]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1086\, Y => 
        \MemorySynchronizer_0/N_1117\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[3]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[3]\, B => 
        \sb_sb_0_Memory_PRDATA[3]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[27]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[27]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[27]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[27]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[23]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[23]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[25]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[23]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[9]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[9]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1[23]\, Y => 
        \MemorySynchronizer_0/N_1082\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_153\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/TimeStampGen/counter[5]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[5]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_41_set_RNIVFGK\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_41_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[19]\, C => 
        \MemorySynchronizer_0/un1_nreset_14_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[19]\);
    
    \STAMP_0/PREADY_0_sqmuxa_2_0_a3\ : CFG4
      generic map(INIT => x"8C0C")

      port map(A => \STAMP_0/apb_spi_finished_Z\, B => 
        \STAMP_0/component_state_Z[3]\, C => 
        \STAMP_0/un13_paddr_i_0\, D => \STAMP_0/un27_paddr_i_0\, 
        Y => \STAMP_0/PREADY_0_sqmuxa_2\);
    
    \MemorySynchronizer_0/SynchStatusReg2[18]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[18]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[18]\);
    
    \STAMP_0/config[11]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[11]\);
    
    \MemorySynchronizer_0/PRDATA[15]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[15]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[15]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_31\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14]\, 
        IPC => OPEN);
    
    \STAMP_0/status_async_cycles_lm_0[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/status_async_cycles_3_sqmuxa\, B => 
        \STAMP_0/status_async_cycles_s[3]\, C => 
        \STAMP_0/status_async_cycles_1_sqmuxa_Z\, Y => 
        \STAMP_0/status_async_cycles_lm[3]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4[9]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[9]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[9]\, C => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[9]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_8\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[8]\, 
        B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_7_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_8_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_8_Z\, 
        CC => NET_CC_CONFIG651, P => NET_CC_CONFIG649, UB => 
        NET_CC_CONFIG650);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_60_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_15\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_60_set_Z\);
    
    \STAMP_0/un1_spi_rx_data_1[19]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[51]\, B => 
        \STAMP_0/dummy_Z[19]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_636\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_26\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[26]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_25_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[6]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_26_Z\, CC
         => NET_CC_CONFIG375, P => NET_CC_CONFIG373, UB => 
        NET_CC_CONFIG374);
    
    \STAMP_0/drdy_flank_detected_dms1\ : SLE
      port map(D => \STAMP_0/stamp0_ready_dms1_c_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/drdy_flank_detected_dms1_1_sqmuxa_1_i_Z\, ALn
         => \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/drdy_flank_detected_dms1_Z\);
    
    AFLSDF_INV_13 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_46_Z\, Y => 
        \AFLSDF_INV_13\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_1_RNIIGV43\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[3]\, 
        B => \MemorySynchronizer_0/un120_in_enable_a_4[2]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[3]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[2]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[0]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[1]\, CC
         => NET_CC_CONFIG1120, P => NET_CC_CONFIG1118, UB => 
        NET_CC_CONFIG1119);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_25\ : 
        CFG4
      generic map(INIT => x"1000")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[14]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[12]\, C => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_10_Z[20]\, 
        D => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_19_Z\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_25_Z\);
    
    \MemorySynchronizer_0/resettimercounter[20]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_13_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[20]\);
    
    \STAMP_0/spi/clk_toggles_lm_0[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/spi/ss_n_buffer_1_sqmuxa\, B => 
        \STAMP_0/spi/clk_toggles_s_Z[5]\, Y => 
        \STAMP_0/spi/clk_toggles_lm[5]\);
    
    \STAMP_0/un5_async_prescaler_count_s_11\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[11]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_10_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_s_11_S\, Y => OPEN, 
        FCO => OPEN, CC => NET_CC_CONFIG513, P => 
        NET_CC_CONFIG511, UB => NET_CC_CONFIG512);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[24]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[24]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[8]\, Y => 
        \MemorySynchronizer_0/N_1067\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_10\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/PLL_ARST_N_net\, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX2_HOLD_N_net\, IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data_1[23]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[55]\, B => 
        \STAMP_0/dummy_Z[23]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_640\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[21]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[21]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[21]\);
    
    \STAMP_0/spi/busy_7_0_0\ : CFG4
      generic map(INIT => x"4EEE")

      port map(A => \STAMP_0/spi/state_Z[0]\, B => 
        \STAMP_0/enable\, C => \STAMP_0/spi/un7_count_NE_i\, D
         => \STAMP_0/spi/un10_count_i\, Y => \STAMP_0/spi/busy_7\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_181\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_16\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/GPD2_ARST_N_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[6]\);
    
    \MemorySynchronizer_0/resynctimercounter[3]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1119\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[3]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[28]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[28]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[4]\, Y => 
        \MemorySynchronizer_0/N_1063\);
    
    \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0\ : CFG4
      generic map(INIT => x"CCCE")

      port map(A => ENABLE_MEMORY_LED_c, B => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, C => 
        \MemorySynchronizer_0/MemorySyncState_Z[4]\, D => 
        \MemorySynchronizer_0/MemorySyncState_Z[1]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0_Z\);
    
    \MemorySynchronizer_0/enableTimestampGen\ : SLE
      port map(D => ENABLE_MEMORY_LED_c, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/enableTimestampGen_Z\);
    
    \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_1_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \STAMP_0/spi_request_for_Z[1]\, B => 
        \STAMP_0/spi_request_for_Z[0]\, C => 
        \STAMP_0/component_state_Z[0]\, D => \STAMP_0/N_331\, Y
         => \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_1\);
    
    \MemorySynchronizer_0/numberofnewavails_RNIVL541_0[0]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[2]\, 
        B => \MemorySynchronizer_0/numberofnewavails_Z[1]\, C => 
        \MemorySynchronizer_0/numberofnewavails_Z[0]\, Y => 
        \MemorySynchronizer_0/N_2313\);
    
    \STAMP_0/component_state_ns_0_i_a3_1_1[0]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \STAMP_0/component_state_Z[0]\, B => 
        \STAMP_0/N_238\, C => \STAMP_0/N_167\, Y => 
        \STAMP_0/component_state_ns_0_i_a3_1_1_Z[0]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_24\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[24]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[24]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_23\, S => 
        \MemorySynchronizer_0/temp_1[24]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_24\, CC => 
        NET_CC_CONFIG271, P => NET_CC_CONFIG269, UB => 
        NET_CC_CONFIG270);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[15]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[15]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[15]\, C => 
        \MemorySynchronizer_0/N_2598\, D => 
        \MemorySynchronizer_0/N_2576\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[15]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_28\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_129\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_7_RNIKP5B7\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[9]\, 
        B => \MemorySynchronizer_0/un120_in_enable_a_4[8]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[9]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[8]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[3]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[4]\, CC
         => NET_CC_CONFIG1129, P => NET_CC_CONFIG1127, UB => 
        NET_CC_CONFIG1128);
    
    \STAMP_0/un1_spi_rx_data_2[1]\ : CFG4
      generic map(INIT => x"D155")

      port map(A => \STAMP_0/un1_spi_rx_data_2_1_0_Z[1]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/dummy_Z[1]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_651\);
    
    \STAMP_0/spi/tx_buffer[12]\ : SLE
      port map(D => \STAMP_0/spi/N_123\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[12]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[23]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[23]\, B => 
        \MemorySynchronizer_0/un104_in_enable_23\, C => 
        \MemorySynchronizer_0/N_2574\, D => 
        \MemorySynchronizer_0/N_2577\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[23]\);
    
    AFLSDF_INV_16 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_16\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_125\ : 
        IP_INTERFACE
      port map(A => \sb_sb_0/Memory_0_intr_or_0_Y\, B => 
        ADLIB_GND0, C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_23\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[23]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_22_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[23]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_23_Z\, 
        CC => NET_CC_CONFIG173, P => NET_CC_CONFIG171, UB => 
        NET_CC_CONFIG172);
    
    \MemorySynchronizer_0/un1_nreset_4_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_41\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_4_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_4_rs_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[30]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[30]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[30]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[2]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[30]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_263\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[12]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[12]\, B => 
        \sb_sb_0_STAMP_PWDATA[12]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[12]\);
    
    \MemorySynchronizer_0/SynchStatusReg[27]\ : SLE
      port map(D => \MemorySynchronizer_0/N_2035_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[27]\);
    
    \STAMP_0/un1_spi_rx_data[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0/N_650\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_5\, C => 
        \STAMP_0/spi_rx_data[0]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[0]\);
    
    \MemorySynchronizer_0/waitingtimercounter[3]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_2_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[3]\);
    
    \MemorySynchronizer_0/resettimercounter_RNIGMCU[8]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_33_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[8]\, C => 
        \MemorySynchronizer_0/un1_nreset_61_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[8]\);
    
    \STAMP_0/un1_component_state_13_i_a3_0_0\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \STAMP_0/spi_request_for_Z[1]\, B => 
        \STAMP_0/spi_busy\, C => \STAMP_0/N_238\, D => 
        \STAMP_0/spi_request_for_Z[0]\, Y => 
        \STAMP_0/un1_component_state_13_i_a3_0_0_Z\);
    
    \STAMP_0/dummy[28]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_16\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[28]\);
    
    \MemorySynchronizer_0/ConfigReg[21]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[21]\);
    
    AFLSDF_INV_25 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_51_Z\, Y => 
        \AFLSDF_INV_25\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_27\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[27]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_26_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[5]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_27_Z\, CC
         => NET_CC_CONFIG378, P => NET_CC_CONFIG376, UB => 
        NET_CC_CONFIG377);
    
    \MemorySynchronizer_0/PRDATA[18]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[18]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[18]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[16]\ : SLE
      port map(D => \STAMP_0_data_frame[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[16]\);
    
    AFLSDF_INV_85 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_61\, Y => 
        \AFLSDF_INV_85\);
    
    \STAMP_0/measurement_dms2[1]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[33]\);
    
    \STAMP_0/spi/count_cry[27]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[27]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[26]\, S => 
        \STAMP_0/spi/count_s[27]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[27]\, CC => NET_CC_CONFIG1006, P
         => NET_CC_CONFIG1004, UB => NET_CC_CONFIG1005);
    
    \STAMP_0/config[19]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[19]\);
    
    \STAMP_0/spi/count_lm_0[25]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[25]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[25]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[28]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[28]\, B => 
        \MemorySynchronizer_0/un104_in_enable_28\, C => 
        \MemorySynchronizer_0/N_2574\, D => 
        \MemorySynchronizer_0/N_2577\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[28]\);
    
    \STAMP_0/delay_counter_lm_0[19]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[19]\, Y => 
        \STAMP_0/delay_counter_lm[19]\);
    
    \STAMP_0/delay_counter_lm_0[13]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[13]\, Y => 
        \STAMP_0/delay_counter_lm[13]\);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_17\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[19]\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[15]\, C => 
        \MemorySynchronizer_0/waitingtimercounter_Z[5]\, D => 
        \MemorySynchronizer_0/waitingtimercounter_Z[2]\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_17_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[23]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_23_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_84\);
    
    \STAMP_0/un1_spi_rx_data_1[17]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[49]\, B => 
        \STAMP_0/dummy_Z[17]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_634\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14[30]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[30]\, 
        B => \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2567\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1222\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_2\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[2]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_1_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[2]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_2_Z\, 
        CC => NET_CC_CONFIG110, P => NET_CC_CONFIG108, UB => 
        NET_CC_CONFIG109);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[14]\ : SLE
      port map(D => \STAMP_0_data_frame[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[14]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[8]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[8]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1[24]\, Y => 
        \MemorySynchronizer_0/N_1083\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_28\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un104_in_enable_28\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[28]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_27_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_28_Z\, CC => 
        NET_CC_CONFIG907, P => NET_CC_CONFIG905, UB => 
        NET_CC_CONFIG906);
    
    \MemorySynchronizer_0/ReadInterrupt_0_sqmuxa_2_i_0_0\ : CFG4
      generic map(INIT => x"FBFA")

      port map(A => \MemorySynchronizer_0/N_2439\, B => 
        \MemorySynchronizer_0/MemorySyncState_Z[1]\, C => 
        \MemorySynchronizer_0/N_191\, D => 
        \MemorySynchronizer_0/SynchStatusReg_2_sqmuxa_1\, Y => 
        \MemorySynchronizer_0/ReadInterrupt_0_sqmuxa_2_i_0_0_Z\);
    
    \STAMP_0/delay_counter_lm_0[6]\ : CFG4
      generic map(INIT => x"FCAC")

      port map(A => \STAMP_0/N_216_i\, B => 
        \STAMP_0/delay_counter_s[6]\, C => 
        \STAMP_0/component_state_RNIFR114_Z[0]\, D => 
        \STAMP_0/apb_spi_finished_0_sqmuxa_1\, Y => 
        \STAMP_0/delay_counter_lm[6]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_162\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \STAMP_0/spi/tx_buffer_RNO[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[7]\, B => 
        \STAMP_0/spi/tx_buffer_Z[6]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_128\);
    
    \MemorySynchronizer_0/N_2539_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_17\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_2539_set_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[12]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_12\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[12]\, 
        C => \MemorySynchronizer_0/N_1521\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[12]\);
    
    \STAMP_0/apb_is_reset_RNIQDSK\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/component_state_Z[2]\, B => 
        sb_sb_0_STAMP_PENABLE, C => \STAMP_0/apb_is_reset_Z\, Y
         => \STAMP_0/N_329\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[20]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[20]\, B => 
        \sb_sb_0_STAMP_PWDATA[20]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[20]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[11]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[11]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[11]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[11]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_9\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[9]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[9]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_8_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_9_Z\, CC => 
        NET_CC_CONFIG850, P => NET_CC_CONFIG848, UB => 
        NET_CC_CONFIG849);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[18]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_18_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_80\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_4\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_35_set_RNIFIDO\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_35_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[14]\, C => 
        \MemorySynchronizer_0/un1_nreset_7_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[14]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_34_set_RNILOBL\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_34_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[29]\, C => 
        \MemorySynchronizer_0/un1_nreset_8_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[29]\);
    
    \STAMP_0/spi/clk_toggles[1]\ : SLE
      port map(D => \STAMP_0/spi/clk_toggles_lm[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB14_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_37_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/clk_toggles_Z[1]\);
    
    \MemorySynchronizer_0/resettimercounter_RNI1S2V[17]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_43_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[17]\, C => 
        \MemorySynchronizer_0/un1_nreset_16_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[17]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_62\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_14\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_15\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_13_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[15]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_14_Z\, CC
         => NET_CC_CONFIG1065, P => NET_CC_CONFIG1063, UB => 
        NET_CC_CONFIG1064);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[4]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[4]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[15]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[15]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_126\ : 
        IP_INTERFACE
      port map(A => STAMP_0_new_avail, B => ADLIB_GND0, C => 
        ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_265\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_36_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[5]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_36\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_22\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_23\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_21_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[23]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_22_Z\, CC
         => NET_CC_CONFIG1089, P => NET_CC_CONFIG1087, UB => 
        NET_CC_CONFIG1088);
    
    \MemorySynchronizer_0/un1_nreset_39_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[26]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_39_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_224\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_22\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[22]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_21_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[22]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_22_Z\, 
        CC => NET_CC_CONFIG170, P => NET_CC_CONFIG168, UB => 
        NET_CC_CONFIG169);
    
    \STAMP_0/component_state_RNIT8HJ[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/spi_busy\, B => 
        \STAMP_0/component_state_Z[1]\, Y => \STAMP_0/N_216_i\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_60_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[6]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_60\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[19]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[19]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1072\, Y => 
        \MemorySynchronizer_0/N_1103\);
    
    \MemorySynchronizer_0/un1_nreset_1_rs_RNIRAIK\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_49_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[1]\, C
         => \MemorySynchronizer_0/un1_nreset_1_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[1]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_RNO_1[5]\ : 
        CFG4
      generic map(INIT => x"AEFF")

      port map(A => \MemorySynchronizer_0/N_2604\, B => 
        \MemorySynchronizer_0/N_140_2\, C => 
        \MemorySynchronizer_0/SynchStatusReg_N_3_mux\, D => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, Y
         => \MemorySynchronizer_0/SynchStatusReg_N_7\);
    
    \MemorySynchronizer_0/un1_nreset_5_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[5]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_5_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_159\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[28]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[28]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[27]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[28]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[28]\, CC
         => NET_CC_CONFIG90, P => NET_CC_CONFIG88, UB => 
        NET_CC_CONFIG89);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[11]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[11]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[10]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[11]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[11]\, CC
         => NET_CC_CONFIG39, P => NET_CC_CONFIG37, UB => 
        NET_CC_CONFIG38);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_155\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \STAMP_0/spi/clk_toggles[3]\ : SLE
      port map(D => \STAMP_0/spi/clk_toggles_lm[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB14_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_37_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/clk_toggles_Z[3]\);
    
    \LED_RECORDING_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => LED_RECORDING_c, E => ADLIB_VCC1, DOUT => 
        \LED_RECORDING_obuf/U0/DOUT1\, EOUT => 
        \LED_RECORDING_obuf/U0/EOUT1\);
    
    \AND2_0_RNIKOS1/U0_RGB1_RGB6\ : RGB_NG
      port map(An => \AND2_0_RNIKOS1/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB6_rgbr_net_1\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[30]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[30]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[29]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[30]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[30]\, CC
         => NET_CC_CONFIG96, P => NET_CC_CONFIG94, UB => 
        NET_CC_CONFIG95);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[6]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[6]\, B => 
        \MemorySynchronizer_0/N_2567\, C => 
        \MemorySynchronizer_0/N_2586\, Y => 
        \MemorySynchronizer_0/N_1254\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[17]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[17]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[17]\, C => 
        \MemorySynchronizer_0/N_2598\, D => 
        \MemorySynchronizer_0/N_2576\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[17]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_54_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_18\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_54_set_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[13]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[13]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[13]\, C => 
        \MemorySynchronizer_0/N_2593\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[13]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[11]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_11_S\, 
        Y => \MemorySynchronizer_0/N_1537\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[29]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[29]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[3]\, Y => 
        \MemorySynchronizer_0/N_1062\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[7]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[7]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[7]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[7]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_1_0[7]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[7]\);
    
    \SCLK_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \SCLK_obuf/U0/EOUT1\, Y => 
        \SCLK_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/waitingtimercounter[6]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_60_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[6]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[4]\, 
        B => \sb_sb_0_STAMP_PWDATA[4]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[4]\);
    
    \STAMP_0/spi/count[22]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[22]\);
    
    \STAMP_0/measurement_dms1[8]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[56]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[31]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[31]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_Z[31]\);
    
    \STAMP_0/spi/count_cry[1]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[1]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_s_389_FCO\, S => 
        \STAMP_0/spi/count_s[1]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[1]\, CC => NET_CC_CONFIG928, P
         => NET_CC_CONFIG926, UB => NET_CC_CONFIG927);
    
    \MemorySynchronizer_0/SynchStatusReg2[22]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[22]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[22]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_0\ : 
        IP_INTERFACE
      port map(A => \sb_sb_0/PREADY_0_iv_i\, B => ADLIB_VCC1, C
         => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net\, IPB
         => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0[30]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[30]\, B => 
        \sb_sb_0_STAMP_PWDATA[30]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[30]\);
    
    \STAMP_0/un1_spi_rx_data_1[20]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[52]\, B => 
        \STAMP_0/dummy_Z[20]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_637\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa_i_1_i_a2\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa_i_1_i_a2_1_Z\, 
        B => \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_271\, D => 
        \MemorySynchronizer_0/N_2569\, Y => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\);
    
    \MemorySynchronizer_0/un1_nreset_52_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[14]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_52_i\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_15\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[15]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_14_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_15_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_15_Z\, 
        CC => NET_CC_CONFIG672, P => NET_CC_CONFIG670, UB => 
        NET_CC_CONFIG671);
    
    \STAMP_0/component_state_RNII1E02[0]\ : CFG4
      generic map(INIT => x"5510")

      port map(A => \STAMP_0/component_state_Z[5]\, B => 
        \STAMP_0/component_state_Z[0]\, C => \STAMP_0/N_168\, D
         => \STAMP_0/N_353\, Y => \STAMP_0/N_263\);
    
    \MemorySynchronizer_0/ConfigReg_RNO[29]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sb_sb_0_STAMP_PWDATA[29]\, B => 
        \MemorySynchronizer_0/APBState_Z[1]\, Y => 
        \MemorySynchronizer_0/N_2305_i\);
    
    \STAMP_0/spi_request_for_RNO[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/spi_dms2_cs_1_sqmuxa_1\, B => 
        \STAMP_0/component_state_Z[3]\, Y => \STAMP_0/N_567_i\);
    
    \stamp0_spi_miso_ibuf/U0/U_IOINFF\ : IOINFF_BYPASS
      port map(A => \stamp0_spi_miso_ibuf/U0/YIN1\, Y => 
        \stamp0_spi_miso_ibuf/U0/YIN\);
    
    \STAMP_0/status_temp_overwrittenVal_9\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/un1_new_avail_0_sqmuxa_1\, B => 
        \STAMP_0_data_frame[13]\, Y => 
        \STAMP_0/status_temp_overwrittenVal_9_Z\);
    
    \MemorySynchronizer_0/resynctimercounter[27]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1095\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[27]\);
    
    \MemorySynchronizer_0/PRDATA[11]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[11]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[11]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[14]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[14]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[14]\);
    
    \STAMP_0/spi/un7_count_NE_17\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \STAMP_0/spi/count_Z[15]\, B => 
        \STAMP_0/spi/count_Z[14]\, C => \STAMP_0/spi/count_Z[13]\, 
        D => \STAMP_0/spi/count_Z[12]\, Y => 
        \STAMP_0/spi/un7_count_NE_17_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO[23]\ : CFG4
      generic map(INIT => x"050D")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_2_0_Z[20]\, 
        B => \MemorySynchronizer_0/N_2321\, C => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, D => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\, 
        Y => \MemorySynchronizer_0/N_2032_i\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[24]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[24]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1067\, Y => 
        \MemorySynchronizer_0/N_1098\);
    
    \STAMP_0/config_RNI6A0E1[31]\ : CFG4
      generic map(INIT => x"FFE0")

      port map(A => MemorySynchronizer_0_dataReadyReset, B => 
        \STAMP_0/config_Z[31]\, C => 
        \STAMP_0/component_state_Z[5]\, D => \STAMP_0/N_329\, Y
         => \STAMP_0/un1_new_avail_0_sqmuxa_1\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[3]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[3]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1[29]\, Y => 
        \MemorySynchronizer_0/N_1088\);
    
    \STAMP_0/un1_spi_rx_data[9]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_659\, C => \STAMP_0/spi_rx_data[9]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[9]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6[7]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[7]\, B => 
        \MemorySynchronizer_0/un104_in_enable_7\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[7]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[11]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[11]\, B => 
        \sb_sb_0_Memory_PRDATA[11]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_60_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_19\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_60_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_65\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resynceventpulldowncounter_RNO[1]\ : 
        CFG3
      generic map(INIT => x"A6")

      port map(A => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[1]\, B
         => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[0]\, C
         => \MemorySynchronizer_0/N_2333\, Y => 
        \MemorySynchronizer_0/N_527_i_i\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[22]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[22]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[22]\, D
         => \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[22]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[28]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[28]\, B => 
        \sb_sb_0_STAMP_PWDATA[28]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[28]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_48\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2]\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/spi/clk_toggles[5]\ : SLE
      port map(D => \STAMP_0/spi/clk_toggles_lm[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB14_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_37_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/clk_toggles_Z[5]\);
    
    \STAMP_0/un1_component_state_17_i_o2_RNO\ : CFG4
      generic map(INIT => x"D0F0")

      port map(A => \STAMP_0/drdy_flank_detected_dms2_Z\, B => 
        \STAMP_0/drdy_flank_detected_dms1_Z\, C => 
        \STAMP_0/component_state_Z[5]\, D => \STAMP_0/N_363\, Y
         => \STAMP_0/N_112_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_156\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/spi/count_cry[28]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[28]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[27]\, S => 
        \STAMP_0/spi/count_s[28]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[28]\, CC => NET_CC_CONFIG1009, P
         => NET_CC_CONFIG1007, UB => NET_CC_CONFIG1008);
    
    \MemorySynchronizer_0/N_2536_set_RNIE1C8\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_2536_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[0]\, C => 
        \MemorySynchronizer_0/un1_nreset_34_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[0]\);
    
    \MemorySynchronizer_0/ConfigReg[12]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[12]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_4[15]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_15_S\, 
        Y => \MemorySynchronizer_0/N_1213\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_49_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_20\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_49_set_Z\);
    
    \STAMP_0/spi/tx_buffer[8]\ : SLE
      port map(D => \STAMP_0/spi/N_127\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[8]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_6\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[6]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[6]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_5_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_6_Z\, CC => 
        NET_CC_CONFIG841, P => NET_CC_CONFIG839, UB => 
        NET_CC_CONFIG840);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_254\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_20\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[20]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_19_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[12]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_20_Z\, CC
         => NET_CC_CONFIG357, P => NET_CC_CONFIG355, UB => 
        NET_CC_CONFIG356);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_198\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14]\, 
        IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data_0[24]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame[24]\, B => 
        \STAMP_0/config_Z[24]\, C => \sb_sb_0_STAMP_PADDR[8]\, Y
         => \STAMP_0/N_607\);
    
    \STAMP_0/delay_counter_lm_0[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_216_i\, B => 
        \STAMP_0/component_state_RNIFR114_Z[0]\, C => 
        \STAMP_0/delay_counter_s[1]\, Y => 
        \STAMP_0/delay_counter_lm[1]\);
    
    \MemorySynchronizer_0/N_2537_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_21\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_2537_set_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter[29]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[29]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_36_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[29]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[24]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_24\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[24]\, 
        C => \MemorySynchronizer_0/N_2418\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[24]\);
    
    \MemorySynchronizer_0/TimeStampReg[5]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[5]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[5]\);
    
    AFLSDF_INV_107 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_48\, Y => 
        \AFLSDF_INV_107\);
    
    \STAMP_0/un1_spi_rx_data_2_1_0[2]\ : CFG4
      generic map(INIT => x"5553")

      port map(A => \STAMP_0_data_frame[2]\, B => 
        \STAMP_0_data_frame[34]\, C => \sb_sb_0_STAMP_PADDR[9]\, 
        D => \sb_sb_0_STAMP_PADDR[7]\, Y => 
        \STAMP_0/un1_spi_rx_data_2_1_0_Z[2]\);
    
    \MemorySynchronizer_0/resynctimercounter[6]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1116\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[6]\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0_1[0]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \MemorySynchronizer_0/N_2553\, B => 
        \MemorySynchronizer_0/MemorySyncState_Z[4]\, C => 
        \MemorySynchronizer_0/N_1482\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa\, Y => 
        \MemorySynchronizer_0/MemorySyncState_ns_0_1_Z[0]\);
    
    AFLSDF_INV_65 : INV_BA
      port map(A => \MemorySynchronizer_0/N_1980_i\, Y => 
        \AFLSDF_INV_65\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_16\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[21]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[28]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28]\, 
        IPC => OPEN);
    
    AFLSDF_INV_43 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_43\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_4\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[4]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_3_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[4]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_4_Z\, 
        CC => NET_CC_CONFIG116, P => NET_CC_CONFIG114, UB => 
        NET_CC_CONFIG115);
    
    \MemorySynchronizer_0/PRDATA[29]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[29]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[29]\);
    
    \STAMP_0/spi/count_cry[7]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[7]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[6]\, S => 
        \STAMP_0/spi/count_s[7]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[7]\, CC => NET_CC_CONFIG946, P
         => NET_CC_CONFIG944, UB => NET_CC_CONFIG945);
    
    \STAMP_0/config[7]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[7]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[0]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[0]\);
    
    AFLSDF_INV_21 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_52_i_i_a2_Z\, 
        Y => \AFLSDF_INV_21\);
    
    \MemorySynchronizer_0/PRDATA[23]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[23]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[23]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[1]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[1]\, 
        B => \sb_sb_0_STAMP_PWDATA[1]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[1]\);
    
    AFLSDF_INV_81 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_81\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_220\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16]\, 
        IPC => OPEN);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB2\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[18]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_18_S\, 
        Y => \MemorySynchronizer_0/N_1509\);
    
    \RXSM_SODS_ibuf/U0/U_IOIN\ : IOIN_IB
      port map(YIN => \RXSM_SODS_ibuf/U0/YIN\, E => ADLIB_GND0, Y
         => RXSM_SODS_c);
    
    \MemorySynchronizer_0/resettimercounter_RNI0A811[13]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_59_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[13]\, C => 
        \MemorySynchronizer_0/un1_nreset_21_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[13]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg_RNI48CK[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[3]\, B => NN_1, 
        Y => \MemorySynchronizer_0/N_1978_i\);
    
    \MemorySynchronizer_0/SynchStatusReg2[6]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[6]\);
    
    \STAMP_0/un1_spi_rx_data_2[15]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_598\, B => \STAMP_0/N_632\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_665\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_53_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_22\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_53_set_Z\);
    
    \STAMP_0/un1_spi_rx_data_2[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_587\, B => \STAMP_0/N_621\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_654\);
    
    
        \MemorySynchronizer_0/SynchStatusReg_2_sqmuxa_1_0_a2_0_a2_RNI2K0M\ : 
        CFG3
      generic map(INIT => x"0E")

      port map(A => \MemorySynchronizer_0/N_2028_i\, B => 
        \MemorySynchronizer_0/SynchStatusReg_2_sqmuxa_1\, C => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, Y => 
        \MemorySynchronizer_0/N_1512\);
    
    \STAMP_0/PRDATA[11]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[11]\);
    
    \MemorySynchronizer_0/ConfigReg[6]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[6]\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_27\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \MemorySynchronizer_0/N_1085\, B => 
        \MemorySynchronizer_0/N_1075\, C => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_21_Z\, D
         => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_7_Z\, 
        Y => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_27_Z\);
    
    \STAMP_0/spi/count[19]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[19]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_RNIC38O1[0]_CC_1\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO1114, CO => OPEN, P(0) => 
        NET_CC_CONFIG1142, P(1) => NET_CC_CONFIG1145, P(2) => 
        NET_CC_CONFIG1148, P(3) => NET_CC_CONFIG1151, P(4) => 
        NET_CC_CONFIG1154, P(5) => NET_CC_CONFIG1157, P(6) => 
        NET_CC_CONFIG1160, P(7) => NET_CC_CONFIG1163, P(8) => 
        ADLIB_VCC1, P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, 
        P(11) => ADLIB_VCC1, UB(0) => NET_CC_CONFIG1143, UB(1)
         => NET_CC_CONFIG1146, UB(2) => NET_CC_CONFIG1149, UB(3)
         => NET_CC_CONFIG1152, UB(4) => NET_CC_CONFIG1155, UB(5)
         => NET_CC_CONFIG1158, UB(6) => NET_CC_CONFIG1161, UB(7)
         => NET_CC_CONFIG1164, UB(8) => ADLIB_VCC1, UB(9) => 
        ADLIB_VCC1, UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, 
        CC(0) => NET_CC_CONFIG1144, CC(1) => NET_CC_CONFIG1147, 
        CC(2) => NET_CC_CONFIG1150, CC(3) => NET_CC_CONFIG1153, 
        CC(4) => NET_CC_CONFIG1156, CC(5) => NET_CC_CONFIG1159, 
        CC(6) => NET_CC_CONFIG1162, CC(7) => NET_CC_CONFIG1165, 
        CC(8) => nc116, CC(9) => nc74, CC(10) => nc133, CC(11)
         => nc420);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_81\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[27]\, B => 
        \MemorySynchronizer_0/un104_in_enable_26\, C => 
        \MemorySynchronizer_0/un104_in_enable_27\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[26]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[12]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[13]\, CC
         => NET_CC_CONFIG577, P => NET_CC_CONFIG575, UB => 
        NET_CC_CONFIG576);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_41\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[19]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_41_Z\);
    
    \MemorySynchronizer_0/un94_in_enable_16\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[31]\, B => 
        \MemorySynchronizer_0/resettimercounter_Z[18]\, C => 
        \MemorySynchronizer_0/resettimercounter_Z[17]\, D => 
        \MemorySynchronizer_0/resettimercounter_Z[16]\, Y => 
        \MemorySynchronizer_0/un94_in_enable_16_Z\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_1\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[1]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_0_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_1_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_1_Z\, CC
         => NET_CC_CONFIG728, P => NET_CC_CONFIG726, UB => 
        NET_CC_CONFIG727);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_11_RNIPSAP7\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[13]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[12]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[13]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[12]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[5]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[6]\, CC
         => NET_CC_CONFIG1135, P => NET_CC_CONFIG1133, UB => 
        NET_CC_CONFIG1134);
    
    \MemorySynchronizer_0/resynceventpulldowncounter[1]\ : SLE
      port map(D => \MemorySynchronizer_0/N_527_i_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[1]\);
    
    \MemorySynchronizer_0/un1_nreset_18_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/N_1979_i\, EN => ADLIB_VCC1, ALn
         => \MemorySynchronizer_0/un1_nreset_18_i\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_18_rs_Z\);
    
    \MemorySynchronizer_0/resynctimercounter[11]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1111\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[11]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_RNO[30]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_30_S\, 
        Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[1]\);
    
    AFLSDF_INV_46 : INV_BA
      port map(A => \MemorySynchronizer_0/N_1979_i\, Y => 
        \AFLSDF_INV_46\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[5]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_5\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[5]\, 
        C => \MemorySynchronizer_0/N_1553\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[5]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10[10]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \sb_sb_0_STAMP_PADDR[9]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \sb_sb_0_STAMP_PADDR[7]\, 
        D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_N_2L1_Z\, Y
         => \MemorySynchronizer_0/N_271\);
    
    \MemorySynchronizer_0/waitingtimercounter[23]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[23]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_25_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[23]\);
    
    \MemorySynchronizer_0/un1_nreset_9_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_49_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_9_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_9_rs_Z\);
    
    \STAMP_0/dummy[27]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_23\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[27]\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_5\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX1_HOLD_N_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[3]\);
    
    \MemorySynchronizer_0/TimeStampGen/un6_enable_3_RNITPHU\ : 
        CFG4
      generic map(INIT => x"0040")

      port map(A => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[1]\, B => 
        \MemorySynchronizer_0/enableTimestampGen_Z\, C => 
        \MemorySynchronizer_0/TimeStampGen/un6_enable_3_Z\, D => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[0]\, Y => 
        \MemorySynchronizer_0/TimeStampGen/countere\);
    
    \MemorySynchronizer_0/un1_nreset_32_rs_RNI895F\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_51_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[2]\, C => 
        \MemorySynchronizer_0/un1_nreset_32_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[2]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[28]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \MemorySynchronizer_0/N_2588\, B => 
        \MemorySynchronizer_0/N_2597\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[28]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[28]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[28]\);
    
    \STAMP_0/spi/tx_buffer[10]\ : SLE
      port map(D => \STAMP_0/spi/N_125\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[10]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[0]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[0]\, B => 
        \sb_sb_0_STAMP_PWDATA[0]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[0]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[9]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_9\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[9]\, 
        C => \MemorySynchronizer_0/N_1533\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[9]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_161\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_100\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[0]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[7]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_134\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \AND2_0_RNIKOS1/U0_RGB1_RGB5\ : RGB_NG
      port map(An => \AND2_0_RNIKOS1/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB5_rgbr_net_1\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO[5]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/g1\, B => 
        \MemorySynchronizer_0/N_4\, C => 
        \MemorySynchronizer_0/g2\, D => 
        \MemorySynchronizer_0/N_2510\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168[3]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[5]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2585\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[5]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[5]\, D => 
        \MemorySynchronizer_0/N_1365\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[5]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_0[28]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \sb_sb_0_STAMP_PADDR[2]\, B => 
        \sb_sb_0_STAMP_PADDR[4]\, C => \sb_sb_0_STAMP_PADDR[5]\, 
        Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_0_Z[28]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_40_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[22]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_40\);
    
    \MemorySynchronizer_0/ConfigReg[13]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[13]\);
    
    \STAMP_0/un1_component_state_17_i_0\ : CFG4
      generic map(INIT => x"EA00")

      port map(A => \STAMP_0/N_364\, B => \STAMP_0/N_248_2\, C
         => \STAMP_0/spi_request_for_Z[0]\, D => \STAMP_0/N_166\, 
        Y => \STAMP_0/N_46\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[4]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_4_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[28]\);
    
    \MemorySynchronizer_0/un94_in_enable_29\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/un94_in_enable_20_Z\, B
         => \MemorySynchronizer_0/un94_in_enable_23_Z\, C => 
        \MemorySynchronizer_0/un94_in_enable_22_Z\, D => 
        \MemorySynchronizer_0/un94_in_enable_21_Z\, Y => 
        \MemorySynchronizer_0/un94_in_enable_29_Z\);
    
    \STAMP_0/measurement_dms1[4]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[52]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_26\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[14]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[14]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[14]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[18]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[14]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10[13]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[13]\, B => 
        \MemorySynchronizer_0/N_2567\, C => 
        \MemorySynchronizer_0/N_2586\, Y => 
        \MemorySynchronizer_0/N_1236\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_3\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[3]\, 
        B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_2_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_3_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_3_Z\, 
        CC => NET_CC_CONFIG636, P => NET_CC_CONFIG634, UB => 
        NET_CC_CONFIG635);
    
    \STAMP_0/delay_counter_lm_0[9]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[9]\, Y => 
        \STAMP_0/delay_counter_lm[9]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[0]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[0]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_60\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[10]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_60_Z\);
    
    \MemorySynchronizer_0/numberofnewavails_RNIVL541[0]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[2]\, 
        B => \MemorySynchronizer_0/numberofnewavails_Z[1]\, C => 
        \MemorySynchronizer_0/numberofnewavails_Z[0]\, Y => 
        \MemorySynchronizer_0/N_2330\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_0\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[0]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[0]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => ADLIB_VCC1, S => OPEN, 
        Y => \MemorySynchronizer_0/temp_1_cry_0_Y\, FCO => 
        \MemorySynchronizer_0/temp_1_cry_0\, CC => 
        NET_CC_CONFIG199, P => NET_CC_CONFIG197, UB => 
        NET_CC_CONFIG198);
    
    \STAMP_0/spi/tx_buffer[2]\ : SLE
      port map(D => \STAMP_0/spi/N_138\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[2]\);
    
    \STAMP_0/measurement_temp[14]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[30]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_53_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[13]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_53\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[14]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[14]\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2564\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1461\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_15\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/NGMUX3_ARST_N_net\, IPB
         => \sb_sb_0/CCC_0/CCC_INST/GPD1_ARST_N_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[5]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_42_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_24\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_42_set_Z\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_3_RNI0UMH4\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[5]\, 
        B => \MemorySynchronizer_0/un120_in_enable_a_4[4]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[5]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[4]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[1]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[2]\, CC
         => NET_CC_CONFIG1123, P => NET_CC_CONFIG1121, UB => 
        NET_CC_CONFIG1122);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[8]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[8]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[8]\, C => 
        \MemorySynchronizer_0/N_2596\, D => 
        \MemorySynchronizer_0/N_2595\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[8]\);
    
    AFLSDF_INV_39 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_48_Z\, Y => 
        \AFLSDF_INV_39\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_51_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_25\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_51_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_177\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_23[10]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_18_0_Z[19]\, B
         => \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[4]\, Y => 
        \MemorySynchronizer_0/N_1182\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[16]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => \MemorySynchronizer_0/N_2597\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[16]\, C => 
        \MemorySynchronizer_0/TimeStampReg_Z[16]\, D => 
        \MemorySynchronizer_0/N_1228\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[16]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_9\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1[0]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => \MemorySynchronizer_0/N_2509\, B => 
        \MemorySynchronizer_0/N_2510\, C => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_a2_0_Z[0]\, 
        D => \MemorySynchronizer_0/N_2326\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168[0]\);
    
    \STAMP_0/dummy[24]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_26\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[24]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[24]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[24]\, B => 
        \sb_sb_0_STAMP_PWDATA[24]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[24]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_0_a0_0\ : 
        CFG2
      generic map(INIT => x"4")

      port map(A => 
        \MemorySynchronizer_0/un1_in_enable_2_0_0_a2_0_Z\, B => 
        \MemorySynchronizer_0/N_2313\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_N_3_mux\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[27]\ : SLE
      port map(D => \STAMP_0_data_frame[59]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[27]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[19]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[19]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[18]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[19]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[19]\, CC
         => NET_CC_CONFIG63, P => NET_CC_CONFIG61, UB => 
        NET_CC_CONFIG62);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_250\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2]\, 
        IPC => OPEN);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_18\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[6]\, 
        B => \MemorySynchronizer_0/un120_in_enable_i_A[7]\, C => 
        \MemorySynchronizer_0/un120_in_enable_i_A[8]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[9]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_18_Z\);
    
    \STAMP_0/spi_tx_data[1]\ : SLE
      port map(D => \STAMP_0/N_297_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[1]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_s_387_CC_1\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO2, CO => CI_TO_CO3, P(0) => 
        NET_CC_CONFIG31, P(1) => NET_CC_CONFIG34, P(2) => 
        NET_CC_CONFIG37, P(3) => NET_CC_CONFIG40, P(4) => 
        NET_CC_CONFIG43, P(5) => NET_CC_CONFIG46, P(6) => 
        NET_CC_CONFIG49, P(7) => NET_CC_CONFIG52, P(8) => 
        NET_CC_CONFIG55, P(9) => NET_CC_CONFIG58, P(10) => 
        NET_CC_CONFIG61, P(11) => NET_CC_CONFIG64, UB(0) => 
        NET_CC_CONFIG32, UB(1) => NET_CC_CONFIG35, UB(2) => 
        NET_CC_CONFIG38, UB(3) => NET_CC_CONFIG41, UB(4) => 
        NET_CC_CONFIG44, UB(5) => NET_CC_CONFIG47, UB(6) => 
        NET_CC_CONFIG50, UB(7) => NET_CC_CONFIG53, UB(8) => 
        NET_CC_CONFIG56, UB(9) => NET_CC_CONFIG59, UB(10) => 
        NET_CC_CONFIG62, UB(11) => NET_CC_CONFIG65, CC(0) => 
        NET_CC_CONFIG33, CC(1) => NET_CC_CONFIG36, CC(2) => 
        NET_CC_CONFIG39, CC(3) => NET_CC_CONFIG42, CC(4) => 
        NET_CC_CONFIG45, CC(5) => NET_CC_CONFIG48, CC(6) => 
        NET_CC_CONFIG51, CC(7) => NET_CC_CONFIG54, CC(8) => 
        NET_CC_CONFIG57, CC(9) => NET_CC_CONFIG60, CC(10) => 
        NET_CC_CONFIG63, CC(11) => NET_CC_CONFIG66);
    
    AFLSDF_INV_37 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_37\, Y => 
        \AFLSDF_INV_37\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_25\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[25]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[25]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_24\, S => 
        \MemorySynchronizer_0/temp_1[25]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_25\, CC => 
        NET_CC_CONFIG274, P => NET_CC_CONFIG272, UB => 
        NET_CC_CONFIG273);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[31]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[31]\, 
        B => \MemorySynchronizer_0/TimeStampReg_Z[31]\, C => 
        \MemorySynchronizer_0/N_2576\, D => 
        \MemorySynchronizer_0/N_1182\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[31]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_RNO[28]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[2]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[28]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[28]\);
    
    \MemorySynchronizer_0/resettimercounter[24]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_9_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[24]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_25[10]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_2567\, C => 
        \MemorySynchronizer_0/N_271\, Y => 
        \MemorySynchronizer_0/N_2581\);
    
    \MemorySynchronizer_0/numberofnewavails_RNI0D491_0[0]\ : CFG4
      generic map(INIT => x"3337")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[0]\, 
        B => \MemorySynchronizer_0/N_140_2\, C => 
        \MemorySynchronizer_0/numberofnewavails_Z[2]\, D => 
        \MemorySynchronizer_0/numberofnewavails_Z[1]\, Y => 
        \MemorySynchronizer_0/N_2310\);
    
    \MemorySynchronizer_0/un1_nreset_1_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[1]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_1_i\);
    
    \STAMP_0/delay_counter[11]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[11]\);
    
    \MemorySynchronizer_0/un1_nreset_38_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_45\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_38_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_38_rs_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[0]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0_Y\, 
        Y => \MemorySynchronizer_0/N_1557\);
    
    \STAMP_0/un1_spi_rx_data_1[9]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[41]\, B => 
        \STAMP_0/dummy_Z[9]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_626\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[24]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[24]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[24]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[24]\);
    
    \MemorySynchronizer_0/waitingtimercounter[9]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_57_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[9]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_183\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0[6]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[6]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[6]\, C => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[6]\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21[6]\);
    
    \STAMP_0/spi/count_lm_0[10]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[10]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[10]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[13]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[13]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[13]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[13]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[13]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1078\, Y => 
        \MemorySynchronizer_0/N_1109\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[7]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[7]\);
    
    \STAMP_0/status_async_cycles_cry[3]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0_data_frame[6]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/status_async_cycles_cry_Z[2]\, S => 
        \STAMP_0/status_async_cycles_s[3]\, Y => OPEN, FCO => 
        \STAMP_0/status_async_cycles_cry_Z[3]\, CC => 
        NET_CC_CONFIG598, P => NET_CC_CONFIG596, UB => 
        NET_CC_CONFIG597);
    
    \STAMP_0/spi/count_s_389_CC_3\ : CC_CONFIG
      port map(CI => CI_TO_CO922, CO => OPEN, P(0) => 
        NET_CC_CONFIG998, P(1) => NET_CC_CONFIG1001, P(2) => 
        NET_CC_CONFIG1004, P(3) => NET_CC_CONFIG1007, P(4) => 
        NET_CC_CONFIG1010, P(5) => NET_CC_CONFIG1013, P(6) => 
        NET_CC_CONFIG1016, P(7) => ADLIB_VCC1, P(8) => ADLIB_VCC1, 
        P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, P(11) => 
        ADLIB_VCC1, UB(0) => NET_CC_CONFIG999, UB(1) => 
        NET_CC_CONFIG1002, UB(2) => NET_CC_CONFIG1005, UB(3) => 
        NET_CC_CONFIG1008, UB(4) => NET_CC_CONFIG1011, UB(5) => 
        NET_CC_CONFIG1014, UB(6) => NET_CC_CONFIG1017, UB(7) => 
        ADLIB_VCC1, UB(8) => ADLIB_VCC1, UB(9) => ADLIB_VCC1, 
        UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, CC(0) => 
        NET_CC_CONFIG1000, CC(1) => NET_CC_CONFIG1003, CC(2) => 
        NET_CC_CONFIG1006, CC(3) => NET_CC_CONFIG1009, CC(4) => 
        NET_CC_CONFIG1012, CC(5) => NET_CC_CONFIG1015, CC(6) => 
        NET_CC_CONFIG1018, CC(7) => nc238, CC(8) => nc167, CC(9)
         => nc84, CC(10) => nc39, CC(11) => nc72);
    
    \MemorySynchronizer_0/un1_nreset_47_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_33\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_47_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_47_rs_Z\);
    
    \MISO_ibuf/U0/U_IOPAD\ : sdf_IOPAD_IN
      port map(PAD => MISO, Y => \MISO_ibuf/U0/YIN1\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[12]\ : SLE
      port map(D => \STAMP_0_data_frame[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[12]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[30]\ : SLE
      port map(D => \STAMP_0_data_frame[62]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[30]\);
    
    \STAMP_0/status_async_cycles[4]\ : SLE
      port map(D => \STAMP_0/status_async_cycles_lm[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/status_async_cycles_1_sqmuxa_1_i_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[7]\);
    
    \STAMP_0/status_dms2_overwrittenVal_RNO\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/un1_new_avail_0_sqmuxa_1\, B => 
        \STAMP_0_data_frame[14]\, Y => \STAMP_0/N_117_i\);
    
    \STAMP_0/component_state_ns_i_a3_0_o2[4]\ : CFG3
      generic map(INIT => x"BF")

      port map(A => \STAMP_0/apb_spi_finished_Z\, B => 
        \STAMP_0/component_state_Z[3]\, C => 
        \STAMP_0/un13_paddr_i_0\, Y => \STAMP_0/N_219\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[22]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[22]\, B => 
        \sb_sb_0_STAMP_PWDATA[22]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[22]\);
    
    \MemorySynchronizer_0/un1_nreset_46_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[18]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_46_i\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_29\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_30\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_28_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[30]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_FCNET1\, 
        CC => NET_CC_CONFIG1110, P => NET_CC_CONFIG1108, UB => 
        NET_CC_CONFIG1109);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[21]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[21]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[21]\, D
         => \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[21]\);
    
    \MemorySynchronizer_0/un1_nreset_19_0_a3_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[28]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_19_i\);
    
    \STAMP_0/spi/tx_buffer_RNO[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[12]\, B => 
        \STAMP_0/spi/tx_buffer_Z[11]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_123\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_269\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_41_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/N_1981_i\, EN => ADLIB_VCC1, ALn
         => \MemorySynchronizer_0/un1_nreset_41_i\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_41_rs_Z\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[20]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[20]\, B => 
        \sb_sb_0_Memory_PRDATA[20]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[20]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_16_0[28]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sb_sb_0_STAMP_PADDR[5]\, B => 
        \sb_sb_0_STAMP_PADDR[2]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_16_0_Z[28]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_13\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[13]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_12_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[13]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_13_Z\, 
        CC => NET_CC_CONFIG143, P => NET_CC_CONFIG141, UB => 
        NET_CC_CONFIG142);
    
    AFLSDF_INV_111 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_59_Z\, Y => 
        \AFLSDF_INV_111\);
    
    \SCLK_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => SCLK_c, E => ADLIB_VCC1, DOUT => 
        \SCLK_obuf/U0/DOUT1\, EOUT => \SCLK_obuf/U0/EOUT1\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[5]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[5]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1[27]\, Y => 
        \MemorySynchronizer_0/N_1086\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[28]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[28]\, B => 
        \sb_sb_0_Memory_PRDATA[28]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[28]\);
    
    \STAMP_0/spi/rx_buffer[3]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[3]\);
    
    \STAMP_0/spi/count_lm_0[18]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[18]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[18]\);
    
    \STAMP_0/config[14]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[14]\);
    
    \STAMP_0/dummy[12]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_27\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[12]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_27\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[27]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[27]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_26\, S => 
        \MemorySynchronizer_0/temp_1[27]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_27\, CC => 
        NET_CC_CONFIG280, P => NET_CC_CONFIG278, UB => 
        NET_CC_CONFIG279);
    
    \STAMP_0/delay_counter_RNIEFPA[20]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \STAMP_0/delay_counter_Z[23]\, B => 
        \STAMP_0/delay_counter_Z[22]\, C => 
        \STAMP_0/delay_counter_Z[21]\, D => 
        \STAMP_0/delay_counter_Z[20]\, Y => 
        \STAMP_0/N_517_i_0_a2_15\);
    
    \RXSM_SODS_ibuf/U0/U_IOPAD\ : sdf_IOPAD_IN
      port map(PAD => RXSM_SODS, Y => \RXSM_SODS_ibuf/U0/YIN1\);
    
    \MemorySynchronizer_0/TimeStampReg[6]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[6]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[6]\);
    
    ip_interface_inst : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ff_to_start_net, C => 
        ADLIB_VCC1, IPA => OPEN, IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/status_async_cycles_s[5]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0_data_frame[8]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/status_async_cycles_cry_Z[4]\, S => 
        \STAMP_0/status_async_cycles_s_Z[5]\, Y => OPEN, FCO => 
        OPEN, CC => NET_CC_CONFIG604, P => NET_CC_CONFIG602, UB
         => NET_CC_CONFIG603);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[5]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_52\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[5]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[5]\, D
         => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[5]\);
    
    \MemorySynchronizer_0/ConfigReg[30]\ : SLE
      port map(D => \MemorySynchronizer_0/N_2306_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/un1_APBState_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[30]\);
    
    \MemorySynchronizer_0/resynctimercounter[29]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1093\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[29]\);
    
    \STAMP_0/un1_component_state_14_i_o2\ : CFG2
      generic map(INIT => x"D")

      port map(A => \STAMP_0/N_110_i\, B => 
        \STAMP_0/config_Z[31]\, Y => \STAMP_0/N_165\);
    
    \MemorySynchronizer_0/un1_nreset_45_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[2]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_45_i\);
    
    \MemorySynchronizer_0/un1_nreset_42_rs_RNIT2TI\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_50_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[24]\, C
         => \MemorySynchronizer_0/un1_nreset_42_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[24]\);
    
    AFLSDF_INV_61 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_43\, Y => 
        \AFLSDF_INV_61\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_227\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23]\, 
        IPC => OPEN);
    
    \STAMP_0/spi/rx_buffer[6]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[6]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_1\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[1]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[1]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_1_Z\, 
        CC => NET_CC_CONFIG107, P => NET_CC_CONFIG105, UB => 
        NET_CC_CONFIG106);
    
    \MemorySynchronizer_0/un104_in_enable_cry_12\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[12]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[12]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_11_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_12_Z\, CC => 
        NET_CC_CONFIG859, P => NET_CC_CONFIG857, UB => 
        NET_CC_CONFIG858);
    
    \MemorySynchronizer_0/TimeStampGen/counter[27]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[27]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[27]\);
    
    \STAMP_0/spi_tx_data[6]\ : SLE
      port map(D => \STAMP_0/N_292_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[6]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_0[15]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[15]\, B => 
        \sb_sb_0_STAMP_PWDATA[15]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_0_Z[15]\);
    
    \STAMP_0/un1_spi_rx_data_2_1_0[1]\ : CFG4
      generic map(INIT => x"5553")

      port map(A => \STAMP_0_data_frame[1]\, B => 
        \STAMP_0_data_frame[33]\, C => \sb_sb_0_STAMP_PADDR[9]\, 
        D => \sb_sb_0_STAMP_PADDR[7]\, Y => 
        \STAMP_0/un1_spi_rx_data_2_1_0_Z[1]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_98\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDIF_net\, IPB
         => OPEN, IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_147\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_18\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_19\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_17_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[19]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_18_Z\, CC
         => NET_CC_CONFIG1077, P => NET_CC_CONFIG1075, UB => 
        NET_CC_CONFIG1076);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[25]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[25]\, B => 
        \sb_sb_0_STAMP_PWDATA[25]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[25]\);
    
    \MemorySynchronizer_0/un1_nreset_29_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_48_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_29_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_29_rs_Z\);
    
    \MemorySynchronizer_0/un1_nreset_26_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[25]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_26_i\);
    
    \MemorySynchronizer_0/numberofnewavails[1]\ : SLE
      port map(D => \MemorySynchronizer_0/ConfigReg_Z[1]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/numberofnewavails_0_sqmuxa\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/numberofnewavails_Z[1]\);
    
    \STAMP_0/PRDATA[17]\ : SLE
      port map(D => \STAMP_0/N_667\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_28\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[17]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_7\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[7]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[7]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_6\, S => 
        \MemorySynchronizer_0/temp_1[7]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_7\, CC => 
        NET_CC_CONFIG220, P => NET_CC_CONFIG218, UB => 
        NET_CC_CONFIG219);
    
    \STAMP_0/un1_spi_rx_data_1[25]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[57]\, B => 
        \STAMP_0/dummy_Z[25]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_642\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_21[10]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[2]\, D => \sb_sb_0_STAMP_PADDR[3]\, 
        Y => \MemorySynchronizer_0/N_2575\);
    
    \STAMP_0/un1_spi_rx_data_1[13]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[45]\, B => 
        \STAMP_0/dummy_Z[13]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_630\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[10]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[10]\);
    
    \ENABLE_MEMORY_LED_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \ENABLE_MEMORY_LED_obuf/U0/DOUT1\, Y => 
        \ENABLE_MEMORY_LED_obuf/U0/DOUT\);
    
    \nCS1_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \nCS1_obuf/U0/EOUT1\, Y => 
        \nCS1_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0[19]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[19]\, B => 
        \sb_sb_0_STAMP_PWDATA[19]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[19]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_13\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[13]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_12_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_13_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_13_Z\, CC
         => NET_CC_CONFIG764, P => NET_CC_CONFIG762, UB => 
        NET_CC_CONFIG763);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6[5]\ : CFG4
      generic map(INIT => x"FFBA")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[5]\, B => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[5]\, C => 
        \MemorySynchronizer_0/N_2574\, D => 
        \MemorySynchronizer_0/N_1123\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[5]\);
    
    AFLSDF_INV_53 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_45\, Y => 
        \AFLSDF_INV_53\);
    
    \STAMP_0/PRDATA[8]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[8]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_128\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_12\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[12]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_11_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[12]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_12_Z\, 
        CC => NET_CC_CONFIG140, P => NET_CC_CONFIG138, UB => 
        NET_CC_CONFIG139);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0_0[1]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[2]\, 
        B => \MemorySynchronizer_0/MemorySyncState_Z[4]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, D
         => \MemorySynchronizer_0/N_2553\, Y => 
        \MemorySynchronizer_0/MemorySyncState_ns_0_0_Z[1]\);
    
    \STAMP_0/component_state_ns_0_1[3]\ : CFG4
      generic map(INIT => x"4C5F")

      port map(A => sb_sb_0_STAMP_PENABLE, B => 
        \STAMP_0/un13_paddr_i_0\, C => 
        \STAMP_0/component_state_Z[2]\, D => 
        \STAMP_0/component_state_Z[3]\, Y => 
        \STAMP_0/component_state_ns_0_1_Z[3]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_46\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[0]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[0]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[0]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[0]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[0]\);
    
    \STAMP_0/delay_counter_lm_0[12]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[12]\, Y => 
        \STAMP_0/delay_counter_lm[12]\);
    
    \MemorySynchronizer_0/un1_nreset_25_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[23]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_25_i\);
    
    \sb_sb_0/CoreAPB3_0/iPSELS_raw_1_0[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \sb_sb_0/STAMP_PADDRS[15]\, B => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx\, Y => 
        \sb_sb_0/CoreAPB3_0/iPSELS_raw_1_0_Z[0]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_RNIKHI89\ : 
        ARI1_CC
      generic map(INIT => x"60990")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_Z\, B
         => \MemorySynchronizer_0/un120_in_enable_i_A[30]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[30]\, D => 
        \MemorySynchronizer_0/un104_in_enable_axb_31\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[14]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_RNIKHI89_FCNET1\, 
        CC => NET_CC_CONFIG1162, P => NET_CC_CONFIG1160, UB => 
        NET_CC_CONFIG1161);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0[27]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[27]\, B => 
        \sb_sb_0_STAMP_PWDATA[27]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[27]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[9]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[9]\);
    
    \STAMP_0/dummy[8]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_29\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[8]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_6\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[3]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[3]\, B => 
        \MemorySynchronizer_0/un104_in_enable_3\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[3]\);
    
    \MemorySynchronizer_0/SynchStatusReg[4]\ : SLE
      port map(D => \MemorySynchronizer_0/SynchStatusReg_168[2]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, 
        EN => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[4]\);
    
    \MemorySynchronizer_0/resettimercounter[16]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_17_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[16]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[30]\, B => 
        \sb_sb_0_Memory_PRDATA[30]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[30]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_26\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[26]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_25_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[26]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_26_Z\, 
        CC => NET_CC_CONFIG182, P => NET_CC_CONFIG180, UB => 
        NET_CC_CONFIG181);
    
    \STAMP_0/un1_component_state_17_i_o2\ : CFG2
      generic map(INIT => x"D")

      port map(A => \STAMP_0/N_112_i\, B => 
        \STAMP_0/config_Z[31]\, Y => \STAMP_0/N_166\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[9]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[9]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[9]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[9]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[9]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[9]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_9[30]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[30]\, 
        B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_16_0_Z[28]\, C
         => \MemorySynchronizer_0/N_1182\, Y => 
        \MemorySynchronizer_0/N_1217\);
    
    \MemorySynchronizer_0/APBState[0]\ : SLE
      port map(D => \MemorySynchronizer_0/APBState_ns[0]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/APBState_Z[0]\);
    
    \MemorySynchronizer_0/TimeStampGen/prescaler_5[4]\ : CFG3
      generic map(INIT => x"12")

      port map(A => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_c4\, B
         => \MemorySynchronizer_0/TimeStampGen/countere\, C => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[4]\, Y => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_5_Z[4]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_9\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[9]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_8_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[23]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_9_Z\, CC
         => NET_CC_CONFIG324, P => NET_CC_CONFIG322, UB => 
        NET_CC_CONFIG323);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO[30]\ : CFG4
      generic map(INIT => x"2AAA")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_152_Z[30]\, B => 
        \MemorySynchronizer_0/N_2588\, C => 
        \MemorySynchronizer_0/APBState_Z[1]\, D => 
        \sb_sb_0_STAMP_PWDATA[29]\, Y => 
        \MemorySynchronizer_0/N_2015_i\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[20]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[20]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[20]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[20]\);
    
    AND2_2 : CFG2
      generic map(INIT => x"8")

      port map(A => sb_sb_0_GPIO_3_M2F, B => ADLIB_VCC1, Y => 
        adc_start_c);
    
    AFLSDF_INV_56 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_56\);
    
    \STAMP_0/spi/un10_count_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \STAMP_0/spi/clk_toggles_Z[5]\, B => 
        \STAMP_0/spi/clk_toggles_Z[0]\, C => 
        \STAMP_0/spi/un10_count_0_a2_0_Z\, D => 
        \STAMP_0/spi/un10_count_0_a2_0_0_Z\, Y => 
        \STAMP_0/spi/un10_count_i\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv[30]\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_30\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[30]\, 
        C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[1]\, D
         => \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, 
        Y => \MemorySynchronizer_0/waitingtimercounter_10[30]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_257\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17]\, 
        IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data_2_1_0[0]\ : CFG4
      generic map(INIT => x"5553")

      port map(A => \STAMP_0_data_frame[0]\, B => 
        \STAMP_0_data_frame[32]\, C => \sb_sb_0_STAMP_PADDR[9]\, 
        D => \sb_sb_0_STAMP_PADDR[7]\, Y => 
        \STAMP_0/un1_spi_rx_data_2_1_0_Z[0]\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_1\ : CFG4
      generic map(INIT => x"000D")

      port map(A => 
        \MemorySynchronizer_0/numberofpendingresyncrequest_Z[0]\, 
        B => \STAMP_0_data_frame[9]\, C => 
        \MemorySynchronizer_0/numberofpendingresyncrequest_Z[2]\, 
        D => 
        \MemorySynchronizer_0/numberofpendingresyncrequest_Z[1]\, 
        Y => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_1_Z\);
    
    \MemorySynchronizer_0/resettimercounter[18]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_15_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[18]\);
    
    \MemorySynchronizer_0/PRDATA[12]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[12]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[12]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0_CC_0\ : 
        CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => CI_TO_CO623, P(0) => 
        ADLIB_GND0, P(1) => NET_CC_CONFIG625, P(2) => 
        NET_CC_CONFIG628, P(3) => NET_CC_CONFIG631, P(4) => 
        NET_CC_CONFIG634, P(5) => NET_CC_CONFIG637, P(6) => 
        NET_CC_CONFIG640, P(7) => NET_CC_CONFIG643, P(8) => 
        NET_CC_CONFIG646, P(9) => NET_CC_CONFIG649, P(10) => 
        NET_CC_CONFIG652, P(11) => NET_CC_CONFIG655, UB(0) => 
        ADLIB_VCC1, UB(1) => NET_CC_CONFIG626, UB(2) => 
        NET_CC_CONFIG629, UB(3) => NET_CC_CONFIG632, UB(4) => 
        NET_CC_CONFIG635, UB(5) => NET_CC_CONFIG638, UB(6) => 
        NET_CC_CONFIG641, UB(7) => NET_CC_CONFIG644, UB(8) => 
        NET_CC_CONFIG647, UB(9) => NET_CC_CONFIG650, UB(10) => 
        NET_CC_CONFIG653, UB(11) => NET_CC_CONFIG656, CC(0) => 
        nc256, CC(1) => NET_CC_CONFIG627, CC(2) => 
        NET_CC_CONFIG630, CC(3) => NET_CC_CONFIG633, CC(4) => 
        NET_CC_CONFIG636, CC(5) => NET_CC_CONFIG639, CC(6) => 
        NET_CC_CONFIG642, CC(7) => NET_CC_CONFIG645, CC(8) => 
        NET_CC_CONFIG648, CC(9) => NET_CC_CONFIG651, CC(10) => 
        NET_CC_CONFIG654, CC(11) => NET_CC_CONFIG657);
    
    \MemorySynchronizer_0/SynchStatusReg_2_sqmuxa_1_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"8")

      port map(A => ENABLE_MEMORY_LED_c, B => 
        \MemorySynchronizer_0/MemorySyncState_Z[2]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_2_sqmuxa_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[18]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[18]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[18]\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[18]\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[18]\);
    
    \STAMP_0/spi/count[16]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[16]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_189\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/spi/count[21]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[21]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_185\ : 
        IP_INTERFACE
      port map(A => MMUART_0_RXD_F2M_c, B => ADLIB_VCC1, C => 
        ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net\, 
        IPC => OPEN);
    
    \STAMP_0/un1_pwdata[11]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[11]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => 
        \STAMP_0/un1_pwdata_Z[11]\);
    
    \STAMP_0/status_async_cycles_cry[1]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0_data_frame[4]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/status_async_cycles_s_388_FCO\, S => 
        \STAMP_0/status_async_cycles_s[1]\, Y => OPEN, FCO => 
        \STAMP_0/status_async_cycles_cry_Z[1]\, CC => 
        NET_CC_CONFIG592, P => NET_CC_CONFIG590, UB => 
        NET_CC_CONFIG591);
    
    \MemorySynchronizer_0/ReadInterrupt_0_sqmuxa_2_i_0_a2_0\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[1]\, 
        B => ENABLE_MEMORY_LED_c, C => 
        \MemorySynchronizer_0/ConfigReg_Z[31]\, D => 
        \MemorySynchronizer_0/end_one_counter_Z[1]\, Y => 
        \MemorySynchronizer_0/N_2439\);
    
    \STAMP_0/spi/un7_count_NE_19\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \STAMP_0/spi/count_Z[7]\, B => 
        \STAMP_0/spi/count_Z[6]\, C => \STAMP_0/spi/count_Z[5]\, 
        D => \STAMP_0/spi/count_Z[4]\, Y => 
        \STAMP_0/spi/un7_count_NE_19_Z\);
    
    \STAMP_0/spi/count[25]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[25]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_13\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[13]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[13]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_12\, S => 
        \MemorySynchronizer_0/temp_1[13]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_13\, CC => 
        NET_CC_CONFIG238, P => NET_CC_CONFIG236, UB => 
        NET_CC_CONFIG237);
    
    \STAMP_0/spi/count_lm_0[26]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[26]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[26]\);
    
    \STAMP_0/component_state[4]\ : SLE
      port map(D => \STAMP_0/component_state_ns[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/component_state_Z[4]\);
    
    \MemorySynchronizer_0/resettimercounter[11]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_3_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[11]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[16]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[16]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1075\, Y => 
        \MemorySynchronizer_0/N_1106\);
    
    \STAMP_0/PRDATA[21]\ : SLE
      port map(D => \STAMP_0/N_671\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_30\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[21]\);
    
    \STAMP_0/spi/ss_n_buffer[0]\ : SLE
      port map(D => \STAMP_0/spi/ss_n_buffer_1_sqmuxa\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/ss_n_buffer_Z[0]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_110\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[2]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[2]\, B => 
        \MemorySynchronizer_0/un104_in_enable_2\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[2]\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_14\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/NGMUX2_ARST_N_net\, IPB
         => \sb_sb_0/CCC_0/CCC_INST/GPD0_ARST_N_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[4]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[28]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_2567\, C => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_2594\);
    
    \sb_sb_0/CCC_0/CCC_INST/INST_CCC_IP\ : CCC

              generic map(INIT => "00" & x"000007FB8000044174000F18C2718C231839DEC0407A04C02501",
         VCOFREQUENCY => 950.000000)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc212, PRDATA(6) => nc205, PRDATA(5) => nc82, 
        PRDATA(4) => nc367, PRDATA(3) => nc145, PRDATA(2) => 
        nc181, PRDATA(1) => nc160, PRDATA(0) => nc57, LOCK => 
        \sb_sb_0/FIC_0_LOCK\, BUSY => OPEN, CLK0 => 
        \sb_sb_0/CCC_0/CCC_INST/CLK0_net\, CLK1 => 
        \sb_sb_0/CCC_0/CCC_INST/CLK1_net\, CLK2 => 
        \sb_sb_0/CCC_0/CCC_INST/CLK2_net\, CLK3 => 
        \sb_sb_0/CCC_0/CCC_INST/CLK3_net\, NGMUX0_SEL => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX0_SEL_net\, NGMUX1_SEL => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX1_SEL_net\, NGMUX2_SEL => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX2_SEL_net\, NGMUX3_SEL => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX3_SEL_net\, NGMUX0_HOLD_N
         => \sb_sb_0/CCC_0/CCC_INST/NGMUX0_HOLD_N_net\, 
        NGMUX1_HOLD_N => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX1_HOLD_N_net\, NGMUX2_HOLD_N
         => \sb_sb_0/CCC_0/CCC_INST/NGMUX2_HOLD_N_net\, 
        NGMUX3_HOLD_N => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX3_HOLD_N_net\, NGMUX0_ARST_N
         => \sb_sb_0/CCC_0/CCC_INST/NGMUX0_ARST_N_net\, 
        NGMUX1_ARST_N => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX1_ARST_N_net\, NGMUX2_ARST_N
         => \sb_sb_0/CCC_0/CCC_INST/NGMUX2_ARST_N_net\, 
        NGMUX3_ARST_N => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX3_ARST_N_net\, PLL_BYPASS_N
         => \sb_sb_0/CCC_0/CCC_INST/PLL_BYPASS_N_net\, PLL_ARST_N
         => \sb_sb_0/CCC_0/CCC_INST/PLL_ARST_N_net\, 
        PLL_POWERDOWN_N => 
        \sb_sb_0/CCC_0/CCC_INST/PLL_POWERDOWN_N_net\, GPD0_ARST_N
         => \sb_sb_0/CCC_0/CCC_INST/GPD0_ARST_N_net\, GPD1_ARST_N
         => \sb_sb_0/CCC_0/CCC_INST/GPD1_ARST_N_net\, GPD2_ARST_N
         => \sb_sb_0/CCC_0/CCC_INST/GPD2_ARST_N_net\, GPD3_ARST_N
         => \sb_sb_0/CCC_0/CCC_INST/GPD3_ARST_N_net\, PRESET_N
         => \sb_sb_0/CCC_0/CCC_INST/PRESET_N_net\, PCLK => 
        \sb_sb_0/CCC_0/CCC_INST/PCLK_net\, PSEL => 
        \sb_sb_0/CCC_0/CCC_INST/PSEL_net\, PENABLE => 
        \sb_sb_0/CCC_0/CCC_INST/PENABLE_net\, PWRITE => 
        \sb_sb_0/CCC_0/CCC_INST/PWRITE_net\, PADDR(7) => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[7]\, PADDR(6) => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[6]\, PADDR(5) => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[5]\, PADDR(4) => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[4]\, PADDR(3) => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[3]\, PADDR(2) => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[2]\, PWDATA(7) => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[7]\, PWDATA(6) => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[6]\, PWDATA(5) => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[5]\, PWDATA(4) => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[4]\, PWDATA(3) => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[3]\, PWDATA(2) => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[2]\, PWDATA(1) => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[1]\, PWDATA(0) => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[0]\, CLK0_PAD => 
        ADLIB_GND0, CLK1_PAD => ADLIB_GND0, CLK2_PAD => 
        ADLIB_GND0, CLK3_PAD => ADLIB_GND0, GL0 => 
        \sb_sb_0/CCC_0/GL0_net\, GL1 => OPEN, GL2 => 
        \sb_sb_0/CCC_0/GL1_net\, GL3 => OPEN, RCOSC_25_50MHZ => 
        \sb_sb_0/FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC\, 
        RCOSC_1MHZ => ADLIB_GND0, XTLOSC => ADLIB_GND0);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[7]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[7]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_8\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[8]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_7_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_8_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_8_Z\, CC
         => NET_CC_CONFIG749, P => NET_CC_CONFIG747, UB => 
        NET_CC_CONFIG748);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_s_30\ : ARI1_CC
      generic map(INIT => x"48F70")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[30]\, B => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, D => 
        \MemorySynchronizer_0/un105_m1_e_0_0\, FCI => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_29_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[30]\, Y
         => OPEN, FCO => OPEN, CC => NET_CC_CONFIG194, P => 
        NET_CC_CONFIG192, UB => NET_CC_CONFIG193);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_0_a2_0_0[22]\ : 
        CFG3
      generic map(INIT => x"DC")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[24]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, C
         => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_0_a2_0_0_Z[22]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_158\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \SCLK_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => SCLK, D => \SCLK_obuf/U0/DOUT\, E => 
        \SCLK_obuf/U0/EOUT\);
    
    \STAMP_0/spi_tx_data[0]\ : SLE
      port map(D => \STAMP_0/N_298_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[0]\);
    
    \STAMP_0/spi/state_RNIDMJE[0]\ : CFG3
      generic map(INIT => x"E0")

      port map(A => \STAMP_0/enable\, B => 
        \STAMP_0/spi/state_Z[0]\, C => debug_led_net_0, Y => 
        \STAMP_0/spi/N_49_i\);
    
    \stamp0_spi_clock_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \stamp0_spi_clock_obuf/U0/EOUT1\, Y => 
        \stamp0_spi_clock_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_30_FCINST1\ : 
        FCEND_BUFF_CC
      port map(FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_FCNET1\, 
        CO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, CC
         => NET_CC_CONFIG390, P => NET_CC_CONFIG388, UB => 
        NET_CC_CONFIG389);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[18]\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \MemorySynchronizer_0/N_2577\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[18]\, C => 
        \MemorySynchronizer_0/un104_in_enable_18\, D => 
        \MemorySynchronizer_0/N_1437\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[18]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[13]\ : SLE
      port map(D => \STAMP_0_data_frame[45]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[13]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[11]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[11]\);
    
    \STAMP_0/PRDATA[16]\ : SLE
      port map(D => \STAMP_0/N_666\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_31\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[16]\);
    
    \MemorySynchronizer_0/un1_nreset_11\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[22]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_11_i\);
    
    \STAMP_0/un1_spi_rx_data_0[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[7]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[7]\, Y
         => \STAMP_0/N_590\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_228\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50]\);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_17\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[17]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[11]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[10]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[3]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_17_Z\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[23]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[23]\);
    
    \STAMP_0/spi_dms1_cs_1_sqmuxa_1_i_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/N_238\, B => \STAMP_0/config_Z[30]\, 
        Y => \STAMP_0/N_363\);
    
    \STAMP_0/delay_counter_cry[11]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[11]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[10]\, S
         => \STAMP_0/delay_counter_s[11]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[11]\, CC => NET_CC_CONFIG428, 
        P => NET_CC_CONFIG426, UB => NET_CC_CONFIG427);
    
    \STAMP_0/status_dms1_overwrittenVal\ : SLE
      port map(D => \STAMP_0/N_116_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_drdy_flank_detected_dms1_0_sqmuxa_1_Z\, ALn
         => \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[12]\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_3\ : IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/PRESET_N_net\, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX1_SEL_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[1]\);
    
    \STAMP_0/un1_spi_rx_data_2[22]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_605\, B => \STAMP_0/N_639\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_672\);
    
    \STAMP_0/spi/count[8]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[8]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[27]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_27\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[23]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[23]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_56_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_32\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_56_set_Z\);
    
    \MemorySynchronizer_0/un1_nreset_3_rs_RNI74OO\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_21_i_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[11]\, C => 
        \MemorySynchronizer_0/un1_nreset_3_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[11]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[26]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[26]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[26]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[26]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_68\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un104_in_enable_cry_7\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[7]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[7]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_6_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_7_Z\, CC => 
        NET_CC_CONFIG844, P => NET_CC_CONFIG842, UB => 
        NET_CC_CONFIG843);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_14[20]\ : 
        CFG2
      generic map(INIT => x"1")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[13]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[16]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_14_Z[20]\);
    
    \STAMP_0/spi/count_s_389_CC_1\ : CC_CONFIG
      port map(CI => CI_TO_CO920, CO => CI_TO_CO921, P(0) => 
        NET_CC_CONFIG926, P(1) => NET_CC_CONFIG929, P(2) => 
        NET_CC_CONFIG932, P(3) => NET_CC_CONFIG935, P(4) => 
        NET_CC_CONFIG938, P(5) => NET_CC_CONFIG941, P(6) => 
        NET_CC_CONFIG944, P(7) => NET_CC_CONFIG947, P(8) => 
        NET_CC_CONFIG950, P(9) => NET_CC_CONFIG953, P(10) => 
        NET_CC_CONFIG956, P(11) => NET_CC_CONFIG959, UB(0) => 
        NET_CC_CONFIG927, UB(1) => NET_CC_CONFIG930, UB(2) => 
        NET_CC_CONFIG933, UB(3) => NET_CC_CONFIG936, UB(4) => 
        NET_CC_CONFIG939, UB(5) => NET_CC_CONFIG942, UB(6) => 
        NET_CC_CONFIG945, UB(7) => NET_CC_CONFIG948, UB(8) => 
        NET_CC_CONFIG951, UB(9) => NET_CC_CONFIG954, UB(10) => 
        NET_CC_CONFIG957, UB(11) => NET_CC_CONFIG960, CC(0) => 
        NET_CC_CONFIG928, CC(1) => NET_CC_CONFIG931, CC(2) => 
        NET_CC_CONFIG934, CC(3) => NET_CC_CONFIG937, CC(4) => 
        NET_CC_CONFIG940, CC(5) => NET_CC_CONFIG943, CC(6) => 
        NET_CC_CONFIG946, CC(7) => NET_CC_CONFIG949, CC(8) => 
        NET_CC_CONFIG952, CC(9) => NET_CC_CONFIG955, CC(10) => 
        NET_CC_CONFIG958, CC(11) => NET_CC_CONFIG961);
    
    \MemorySynchronizer_0/un104_in_enable_cry_21\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[21]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[21]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_20_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_21_Z\, CC => 
        NET_CC_CONFIG886, P => NET_CC_CONFIG884, UB => 
        NET_CC_CONFIG885);
    
    \MemorySynchronizer_0/end_one_counter[1]\ : SLE
      port map(D => \MemorySynchronizer_0/N_2030_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => ADLIB_VCC1, ADn => ADLIB_VCC1, SLn => 
        ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/end_one_counter_Z[1]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_57_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_33\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_57_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_186\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[14]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[3]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[14]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[14]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_1\ : 
        CFG3
      generic map(INIT => x"02")

      port map(A => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, B
         => \MemorySynchronizer_0/N_2604\, C => 
        \MemorySynchronizer_0/un1_enabletimestampgen2_2_sn\, Y
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_1_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_284\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11]\, 
        IPC => OPEN);
    
    \STAMP_0/spi/count[13]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[13]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[25]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[25]\);
    
    \STAMP_0/un1_spi_rx_data_1[10]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[42]\, B => 
        \STAMP_0/dummy_Z[10]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_627\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0_0_0[4]\ : CFG4
      generic map(INIT => x"22F2")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[1]\, 
        B => \MemorySynchronizer_0/end_one_counter_Z[1]\, C => 
        \MemorySynchronizer_0/N_140_2\, D => 
        \MemorySynchronizer_0/MemorySyncState_ns_0_0_0_1_Z[4]\, Y
         => \MemorySynchronizer_0/MemorySyncState_ns[4]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_57_i_i_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[9]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_57_i_i_a2_Z\);
    
    \MemorySynchronizer_0/un1_nreset_10_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[23]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_10_i\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_6\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[6]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_5_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_6_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_6_Z\, CC
         => NET_CC_CONFIG743, P => NET_CC_CONFIG741, UB => 
        NET_CC_CONFIG742);
    
    \STAMP_0/un1_spi_rx_data_0[21]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[21]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[21]\, Y
         => \STAMP_0/N_604\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[13]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[13]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[12]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[13]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[13]\, CC
         => NET_CC_CONFIG45, P => NET_CC_CONFIG43, UB => 
        NET_CC_CONFIG44);
    
    \MemorySynchronizer_0/SynchStatusReg2_RNO[6]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \MemorySynchronizer_0/temp_1_cry_0_Y\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[6]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[6]\);
    
    \MemorySynchronizer_0/un1_nreset_61\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[8]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_61_i\);
    
    \STAMP_0/PRDATA[3]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[3]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[28]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_28\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[28]\, 
        C => \MemorySynchronizer_0/N_1474\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[28]\);
    
    \STAMP_0/spi/count_0_sqmuxa_0_a2\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/enable\, B => 
        \STAMP_0/spi/state_Z[0]\, C => debug_led_net_0, Y => 
        \STAMP_0/spi/count_0_sqmuxa\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_s_387_CC_0\ : 
        CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => CI_TO_CO2, P(0) => 
        ADLIB_VCC1, P(1) => ADLIB_VCC1, P(2) => ADLIB_GND0, P(3)
         => NET_CC_CONFIG4, P(4) => NET_CC_CONFIG7, P(5) => 
        NET_CC_CONFIG10, P(6) => NET_CC_CONFIG13, P(7) => 
        NET_CC_CONFIG16, P(8) => NET_CC_CONFIG19, P(9) => 
        NET_CC_CONFIG22, P(10) => NET_CC_CONFIG25, P(11) => 
        NET_CC_CONFIG28, UB(0) => ADLIB_VCC1, UB(1) => ADLIB_VCC1, 
        UB(2) => ADLIB_GND0, UB(3) => NET_CC_CONFIG5, UB(4) => 
        NET_CC_CONFIG8, UB(5) => NET_CC_CONFIG11, UB(6) => 
        NET_CC_CONFIG14, UB(7) => NET_CC_CONFIG17, UB(8) => 
        NET_CC_CONFIG20, UB(9) => NET_CC_CONFIG23, UB(10) => 
        NET_CC_CONFIG26, UB(11) => NET_CC_CONFIG29, CC(0) => 
        nc430, CC(1) => nc349, CC(2) => nc156, CC(3) => 
        NET_CC_CONFIG6, CC(4) => NET_CC_CONFIG9, CC(5) => 
        NET_CC_CONFIG12, CC(6) => NET_CC_CONFIG15, CC(7) => 
        NET_CC_CONFIG18, CC(8) => NET_CC_CONFIG21, CC(9) => 
        NET_CC_CONFIG24, CC(10) => NET_CC_CONFIG27, CC(11) => 
        NET_CC_CONFIG30);
    
    \MemorySynchronizer_0/resynceventpulldowncounter_RNO[0]\ : 
        CFG2
      generic map(INIT => x"9")

      port map(A => \MemorySynchronizer_0/N_2333\, B => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[0]\, Y
         => \MemorySynchronizer_0/N_1158_i_i\);
    
    \STAMP_0/dummy[31]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[31]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_34\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[31]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_RNO[16]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \MemorySynchronizer_0/temp_1_cry_0_Y\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[16]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[16]\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_i_0_i_a2_0_0[3]\ : 
        CFG4
      generic map(INIT => x"00FE")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[0]\, 
        B => \MemorySynchronizer_0/numberofnewavails_Z[1]\, C => 
        \MemorySynchronizer_0/numberofnewavails_Z[2]\, D => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/un1_in_enable_2_0_0_a2_0_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[12]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[12]\, B => 
        \sb_sb_0_STAMP_PWDATA[12]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[12]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_21[20]\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[30]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[8]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[6]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[1]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_21_Z[20]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[7]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[7]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[7]\, C => 
        \MemorySynchronizer_0/N_2576\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_1_0[7]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_0_a1\ : 
        CFG4
      generic map(INIT => x"2000")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a1_0_0_Z\, 
        B => \sb_sb_0_STAMP_PADDR[5]\, C => 
        \MemorySynchronizer_0/N_271\, D => 
        \MemorySynchronizer_0/N_2567\, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_0_a1_Z\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[11]\ : SLE
      port map(D => \STAMP_0_data_frame[43]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[11]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[15]\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \MemorySynchronizer_0/N_2577\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[15]\, C => 
        \MemorySynchronizer_0/un104_in_enable_15\, D => 
        \MemorySynchronizer_0/N_1453\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[15]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[5]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[5]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[5]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[5]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_163\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA[20]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[20]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[20]\);
    
    \MemorySynchronizer_0/resynctimercounter[7]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1115\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[7]\);
    
    \MemorySynchronizer_0/resynctimercounter[14]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1108\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[14]\);
    
    \STAMP_0/spi_request_for_2_sqmuxa_0_a3\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \STAMP_0/config_Z[30]\, B => 
        \STAMP_0/drdy_flank_detected_temp_Z\, C => 
        \STAMP_0/N_333\, D => \STAMP_0/N_158\, Y => 
        \STAMP_0/spi_request_for_2_sqmuxa\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[12]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[12]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[12]\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[12]\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[12]\);
    
    \STAMP_0/async_state[0]\ : SLE
      port map(D => \STAMP_0/N_90_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/async_state_Z[0]\);
    
    \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1_0_a2\ : 
        CFG4
      generic map(INIT => x"001F")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa\, B => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, C => 
        ENABLE_MEMORY_LED_c, D => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, Y => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\);
    
    \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa_i_0_i_a2_1\ : 
        CFG4
      generic map(INIT => x"0080")

      port map(A => \MemorySynchronizer_0/APBState_Z[1]\, B => 
        \sb_sb_0_STAMP_PADDR[2]\, C => \sb_sb_0_STAMP_PADDR[3]\, 
        D => \sb_sb_0_STAMP_PADDR[6]\, Y => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa_i_0_i_a2_1_Z\);
    
    \STAMP_0/component_state_RNI0A1I[4]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \STAMP_0/component_state_Z[3]\, B => 
        \STAMP_0/component_state_Z[4]\, C => 
        \STAMP_0/component_state_Z[2]\, Y => \STAMP_0/N_163\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[6]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_6\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[6]\, 
        C => \MemorySynchronizer_0/N_1541\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[6]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[29]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[29]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[29]\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[29]\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[29]\);
    
    AFLSDF_INV_34 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_34\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_17\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[17]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_16_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_17_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_17_Z\, CC
         => NET_CC_CONFIG776, P => NET_CC_CONFIG774, UB => 
        NET_CC_CONFIG775);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[9]\ : SLE
      port map(D => \STAMP_0_data_frame[41]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[9]\);
    
    \STAMP_0/spi/count_lm_0[29]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[29]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[29]\);
    
    \STAMP_0/spi_request_for_2_sqmuxa_0_o2_RNI8RIC1\ : CFG4
      generic map(INIT => x"A080")

      port map(A => \STAMP_0/config_Z[30]\, B => 
        \STAMP_0/drdy_flank_detected_temp_Z\, C => 
        \STAMP_0/N_333\, D => \STAMP_0/N_158\, Y => 
        \STAMP_0/N_361\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_258\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg2[19]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[19]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[19]\);
    
    \STAMP_0/dummy[4]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_35\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[4]\);
    
    \STAMP_0/PREADY\ : SLE
      port map(D => \STAMP_0/PREADY_0_sqmuxa_2\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_PREADY_0_sqmuxa_3_0_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => sb_sb_0_STAMP_PREADY);
    
    \MMUART_0_RXD_F2M_ibuf/U0/U_IOIN\ : IOIN_IB
      port map(YIN => \MMUART_0_RXD_F2M_ibuf/U0/YIN\, E => 
        ADLIB_GND0, Y => MMUART_0_RXD_F2M_c);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_20\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[20]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_19_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[20]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_20_Z\, 
        CC => NET_CC_CONFIG164, P => NET_CC_CONFIG162, UB => 
        NET_CC_CONFIG163);
    
    \STAMP_0/async_prescaler_count[1]\ : SLE
      port map(D => \STAMP_0/un5_async_prescaler_count_cry_1_S\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[1]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[8]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[8]\);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.un151_in_enablelto30_17\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/temp_1[21]\, B => 
        \MemorySynchronizer_0/temp_1[22]\, C => 
        \MemorySynchronizer_0/temp_1[23]\, D => 
        \MemorySynchronizer_0/temp_1[24]\, Y => 
        \MemorySynchronizer_0/un151_in_enablelto30_17\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_9\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[9]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[9]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_8\, S => 
        \MemorySynchronizer_0/temp_1[9]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_9\, CC => 
        NET_CC_CONFIG226, P => NET_CC_CONFIG224, UB => 
        NET_CC_CONFIG225);
    
    \RXSM_SOE_ibuf/U0/U_IOPAD\ : sdf_IOPAD_IN
      port map(PAD => RXSM_SOE, Y => \RXSM_SOE_ibuf/U0/YIN1\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[10]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[4]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[10]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[10]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[15]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[4]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[15]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[15]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_18[20]\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[22]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[17]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[15]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[7]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_18_Z[20]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_19\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[19]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[19]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_18_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_19_Z\, CC => 
        NET_CC_CONFIG880, P => NET_CC_CONFIG878, UB => 
        NET_CC_CONFIG879);
    
    \LED_RECORDING_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \LED_RECORDING_obuf/U0/EOUT1\, Y => 
        \LED_RECORDING_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[23]\ : SLE
      port map(D => \STAMP_0_data_frame[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[23]\);
    
    \MemorySynchronizer_0/resettimercounter[6]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[6]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_49_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[6]\);
    
    \MemorySynchronizer_0/un1_nreset_7\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[14]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_7_i\);
    
    \STAMP_0/spi/clk_toggles_cry[2]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/spi/clk_toggles_Z[2]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/spi/clk_toggles_cry_Z[1]\, S
         => \STAMP_0/spi/clk_toggles_s[2]\, Y => OPEN, FCO => 
        \STAMP_0/spi/clk_toggles_cry_Z[2]\, CC => 
        NET_CC_CONFIG613, P => NET_CC_CONFIG611, UB => 
        NET_CC_CONFIG612);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_83\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[26]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[26]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_96\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CRSF_net\, IPB
         => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_32_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[20]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_32\);
    
    \MemorySynchronizer_0/MemorySyncState_RNI5C001[5]\ : CFG4
      generic map(INIT => x"BAFA")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[5]\, 
        B => STAMP_0_new_avail, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, Y
         => \MemorySynchronizer_0/g2_0_0\);
    
    \MemorySynchronizer_0/resynctimercounter[10]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1112\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[10]\);
    
    \STAMP_0/apb_spi_finished\ : SLE
      port map(D => \STAMP_0/un1_apb_spi_finished_1_f0_Z\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN
         => debug_led_net_0, ALn => ADLIB_VCC1, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \STAMP_0/apb_spi_finished_Z\);
    
    \STAMP_0/spi/count_lm_0[11]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[11]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[11]\);
    
    AFLSDF_INV_19 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_60_Z\, Y => 
        \AFLSDF_INV_19\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[9]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[9]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[8]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[9]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[9]\, CC
         => NET_CC_CONFIG33, P => NET_CC_CONFIG31, UB => 
        NET_CC_CONFIG32);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_60_set_RNIND1O\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_60_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[10]\, C => 
        \MemorySynchronizer_0/un1_nreset_23_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[10]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_5_RNIMBEU5\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[7]\, 
        B => \MemorySynchronizer_0/un120_in_enable_a_4[6]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[7]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[6]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[2]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[3]\, CC
         => NET_CC_CONFIG1126, P => NET_CC_CONFIG1124, UB => 
        NET_CC_CONFIG1125);
    
    \MemorySynchronizer_0/waitingtimercounter_RNIH9PT[10]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_2534_set_Z\, B => 
        \MemorySynchronizer_0/waitingtimercounterrs[10]\, C => 
        \MemorySynchronizer_0/un1_nreset_56_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[10]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[25]\ : SLE
      port map(D => \STAMP_0_data_frame[57]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[25]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_N_2L1\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \sb_sb_0_STAMP_PADDR[1]\, B => 
        \sb_sb_0_STAMP_PADDR[11]\, C => \sb_sb_0_STAMP_PADDR[10]\, 
        D => \sb_sb_0_STAMP_PADDR[0]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_N_2L1_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_280\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7]\, 
        IPC => OPEN);
    
    AFLSDF_INV_17 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_32_i_i_a2_Z\, 
        Y => \AFLSDF_INV_17\);
    
    \STAMP_0/request_resync_1_sqmuxa_2_i_0\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/request_resync_1_sqmuxa_1_Z\, B => 
        \STAMP_0/request_resync_0_sqmuxa\, Y => \STAMP_0/N_152\);
    
    \stamp0_spi_dms2_cs_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \stamp0_spi_dms2_cs_obuf/U0/EOUT1\, Y => 
        \stamp0_spi_dms2_cs_obuf/U0/EOUT\);
    
    \STAMP_0/delay_counter[21]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[21]\);
    
    \STAMP_0/PRDATA[27]\ : SLE
      port map(D => \STAMP_0/N_677\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_36\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[27]\);
    
    CFG0_GND_INST : CFG0
      generic map(INIT => "0")

      port map(Y => CFG0_GND_INST_NET);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_10_RNIF76L7\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[11]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[10]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[11]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[10]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[4]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[5]\, CC
         => NET_CC_CONFIG1132, P => NET_CC_CONFIG1130, UB => 
        NET_CC_CONFIG1131);
    
    \MemorySynchronizer_0/numberofpendingresyncrequest[0]\ : SLE
      port map(D => \MemorySynchronizer_0/ConfigReg_Z[4]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN
         => \MemorySynchronizer_0/numberofnewavails_0_sqmuxa\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/numberofpendingresyncrequest_Z[0]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[19]\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \MemorySynchronizer_0/N_2577\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[19]\, C => 
        \MemorySynchronizer_0/un104_in_enable_19\, D => 
        \MemorySynchronizer_0/N_1342\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[19]\);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.un151_in_enablelto30_23\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => 
        \MemorySynchronizer_0/un151_in_enablelto30_14\, B => 
        \MemorySynchronizer_0/un151_in_enablelto30_15\, C => 
        \MemorySynchronizer_0/un151_in_enablelto30_16\, D => 
        \MemorySynchronizer_0/un151_in_enablelto30_17\, Y => 
        \MemorySynchronizer_0/un151_in_enablelto30_23\);
    
    \STAMP_0/delay_counter_lm_0[24]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[24]\, Y => 
        \STAMP_0/delay_counter_lm[24]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_37_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_37\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_37_set_Z\);
    
    \STAMP_0/un1_component_state_9_i_o2_0_RNINUR01\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \STAMP_0/component_state_Z[2]\, B => 
        \STAMP_0/component_state_Z[4]\, C => \STAMP_0/N_160\, D
         => \STAMP_0/component_state_Z[3]\, Y => \STAMP_0/N_168\);
    
    \STAMP_0/spi_tx_data[11]\ : SLE
      port map(D => \STAMP_0/un1_pwdata_Z[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[11]\);
    
    \STAMP_0/delay_counter[17]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[17]\);
    
    \STAMP_0/component_state_ns_0_i_0_0[0]\ : CFG4
      generic map(INIT => x"A0E0")

      port map(A => \STAMP_0/component_state_ns_0_i_0_tz_Z[0]\, B
         => \STAMP_0/component_state_Z[0]\, C => \STAMP_0/N_167\, 
        D => \STAMP_0/N_331\, Y => 
        \STAMP_0/component_state_ns_0_i_0_0_Z[0]\);
    
    \MemorySynchronizer_0/un1_nreset_40_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_31\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_40_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_40_rs_Z\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a1_Z\, 
        B => \MemorySynchronizer_0/N_140_2\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_4_Z\, 
        D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a0_1_Z\, 
        Y => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[30]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[30]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[30]\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB14\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => OPEN, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB14_rgbr_net_1\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_28\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_16_Z\, B => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_17_Z\, C => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_18_Z\, D => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_19_Z\, Y => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_28_Z\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_69\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[25]\, B => 
        \MemorySynchronizer_0/un104_in_enable_24\, C => 
        \MemorySynchronizer_0/un104_in_enable_25\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[24]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[11]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[12]\, CC
         => NET_CC_CONFIG574, P => NET_CC_CONFIG572, UB => 
        NET_CC_CONFIG573);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_24\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[24]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_23_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_24_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_24_Z\, CC
         => NET_CC_CONFIG797, P => NET_CC_CONFIG795, UB => 
        NET_CC_CONFIG796);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_22\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[22]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_21_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_22_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_22_Z\, CC
         => NET_CC_CONFIG791, P => NET_CC_CONFIG789, UB => 
        NET_CC_CONFIG790);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_17[20]\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[29]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[27]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[20]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[9]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_17_Z[20]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_29\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[29]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_28_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[29]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_29_Z\, 
        CC => NET_CC_CONFIG191, P => NET_CC_CONFIG189, UB => 
        NET_CC_CONFIG190);
    
    \STAMP_0/spi/count_cry[25]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[25]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[24]\, S => 
        \STAMP_0/spi/count_s[25]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[25]\, CC => NET_CC_CONFIG1000, P
         => NET_CC_CONFIG998, UB => NET_CC_CONFIG999);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[21]\ : SLE
      port map(D => \STAMP_0_data_frame[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[21]\);
    
    \STAMP_0/un1_spi_rx_data[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0/N_652\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_5\, C => 
        \STAMP_0/spi_rx_data[2]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[2]\);
    
    \MemorySynchronizer_0/SynchStatusReg_152[30]\ : CFG4
      generic map(INIT => x"F9F8")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_152_ss0_i_0\, B => 
        \MemorySynchronizer_0/SynchStatusReg_152_sm0\, C => 
        \MemorySynchronizer_0/SynchStatusReg_Z[30]\, D => 
        \MemorySynchronizer_0/end_one_counter_Z[1]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_152_Z[30]\);
    
    \MemorySynchronizer_0/resettimercounter_2_sqmuxa_0_a2\ : CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa\, C => 
        ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\);
    
    \MemorySynchronizer_0/APBState_ns_1_0_.m3_0_a3_0_a2\ : CFG3
      generic map(INIT => x"02")

      port map(A => sb_sb_0_Memory_PSELx, B => 
        \MemorySynchronizer_0/N_301\, C => sb_sb_0_STAMP_PWRITE, 
        Y => \MemorySynchronizer_0/APBState_ns[0]\);
    
    \MemorySynchronizer_0/resynctimercounter[9]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1113\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[9]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0[28]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \sb_sb_0_STAMP_PADDR[2]\, B => 
        \sb_sb_0_STAMP_PADDR[4]\, C => \sb_sb_0_STAMP_PADDR[5]\, 
        Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_Z[28]\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_17\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_4_S\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_5_S\, 
        C => \MemorySynchronizer_0/un5_resettimercounter_cry_6_S\, 
        D => \MemorySynchronizer_0/un5_resettimercounter_cry_7_S\, 
        Y => \MemorySynchronizer_0/un6_in_enable_0_a3_17_Z\);
    
    \STAMP_0/measurement_dms2[3]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[35]\);
    
    \MemorySynchronizer_0/waitingtimercounter[19]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[19]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbl_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_40_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[19]\);
    
    \MemorySynchronizer_0/resynceventpulldowncounter[2]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1052_i_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[2]\);
    
    \STAMP_0/un1_spi_rx_data_0[12]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[12]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[12]\, Y
         => \STAMP_0/N_595\);
    
    \stamp0_spi_dms1_cs_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => stamp0_spi_dms1_cs_c, E => ADLIB_VCC1, DOUT
         => \stamp0_spi_dms1_cs_obuf/U0/DOUT1\, EOUT => 
        \stamp0_spi_dms1_cs_obuf/U0/EOUT1\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_169\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[2]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[2]\);
    
    \MemorySynchronizer_0/un1_nreset_58_0_a3_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[8]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_58_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_165\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[15]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[15]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[17]\, Y
         => \MemorySynchronizer_0/N_1076\);
    
    \MemorySynchronizer_0/un1_nreset_43_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_39\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_43_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_43_rs_Z\);
    
    \STAMP_0/dummy[22]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_38\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[22]\);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_28\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_22_Z\, B => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_21_Z\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_20_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_19_Z\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\);
    
    \STAMP_0/un1_spi_rx_data[11]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_661\, C => \STAMP_0/spi_rx_data[11]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[11]\);
    
    \STAMP_0/delay_counter_lm_0[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[2]\, Y => 
        \STAMP_0/delay_counter_lm[2]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_197\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_55_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[11]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_55_i\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_48_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_39\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_48_set_Z\);
    
    \STAMP_0/component_state_RNIL8S97[0]\ : CFG4
      generic map(INIT => x"1113")

      port map(A => \STAMP_0/N_238\, B => \STAMP_0/N_263\, C => 
        \STAMP_0/N_353\, D => \STAMP_0/N_168\, Y => 
        \STAMP_0/N_118_i\);
    
    \MemorySynchronizer_0/end_one_counter_RNO[1]\ : CFG3
      generic map(INIT => x"98")

      port map(A => \MemorySynchronizer_0/end_one_counter_Z[1]\, 
        B => \MemorySynchronizer_0/N_2337\, C => 
        \MemorySynchronizer_0/end_one_counter_Z[0]\, Y => 
        \MemorySynchronizer_0/N_2030_i\);
    
    \debug_led_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => debug_led, D => \debug_led_obuf/U0/DOUT\, E
         => \debug_led_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/N_1981_i_set_RNIA84F\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_1981_i_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[12]\, C => 
        \MemorySynchronizer_0/un1_nreset_41_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[12]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_0_a2_0\ : 
        CFG2
      generic map(INIT => x"1")

      port map(A => \sb_sb_0_STAMP_PADDR[4]\, B => 
        \sb_sb_0_STAMP_PADDR[2]\, Y => 
        \MemorySynchronizer_0/N_2569\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[29]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[29]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[29]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_0_CC_1\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO195, CO => CI_TO_CO196, P(0) => 
        NET_CC_CONFIG227, P(1) => NET_CC_CONFIG230, P(2) => 
        NET_CC_CONFIG233, P(3) => NET_CC_CONFIG236, P(4) => 
        NET_CC_CONFIG239, P(5) => NET_CC_CONFIG242, P(6) => 
        NET_CC_CONFIG245, P(7) => NET_CC_CONFIG248, P(8) => 
        NET_CC_CONFIG251, P(9) => NET_CC_CONFIG254, P(10) => 
        NET_CC_CONFIG257, P(11) => NET_CC_CONFIG260, UB(0) => 
        NET_CC_CONFIG228, UB(1) => NET_CC_CONFIG231, UB(2) => 
        NET_CC_CONFIG234, UB(3) => NET_CC_CONFIG237, UB(4) => 
        NET_CC_CONFIG240, UB(5) => NET_CC_CONFIG243, UB(6) => 
        NET_CC_CONFIG246, UB(7) => NET_CC_CONFIG249, UB(8) => 
        NET_CC_CONFIG252, UB(9) => NET_CC_CONFIG255, UB(10) => 
        NET_CC_CONFIG258, UB(11) => NET_CC_CONFIG261, CC(0) => 
        NET_CC_CONFIG229, CC(1) => NET_CC_CONFIG232, CC(2) => 
        NET_CC_CONFIG235, CC(3) => NET_CC_CONFIG238, CC(4) => 
        NET_CC_CONFIG241, CC(5) => NET_CC_CONFIG244, CC(6) => 
        NET_CC_CONFIG247, CC(7) => NET_CC_CONFIG250, CC(8) => 
        NET_CC_CONFIG253, CC(9) => NET_CC_CONFIG256, CC(10) => 
        NET_CC_CONFIG259, CC(11) => NET_CC_CONFIG262);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_37\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20]\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/spi_temp_cs_13_iv_i\ : CFG3
      generic map(INIT => x"13")

      port map(A => \STAMP_0/component_state_Z[3]\, B => 
        \STAMP_0/spi_request_for_2_sqmuxa\, C => 
        \sb_sb_0_STAMP_PADDR[6]\, Y => 
        \STAMP_0/spi_temp_cs_13_iv_i_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[11]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[11]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[11]\, D
         => \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[11]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[3]\ : SLE
      port map(D => \MemorySynchronizer_0/temp_1[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[3]\);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.un151_in_enablelto30_14\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/temp_1[9]\, B => 
        \MemorySynchronizer_0/temp_1[10]\, C => 
        \MemorySynchronizer_0/temp_1[11]\, D => 
        \MemorySynchronizer_0/temp_1[12]\, Y => 
        \MemorySynchronizer_0/un151_in_enablelto30_14\);
    
    \resetn_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \resetn_obuf/U0/DOUT1\, Y => 
        \resetn_obuf/U0/DOUT\);
    
    AFLSDF_INV_72 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_47_i_i_a2_Z\, 
        Y => \AFLSDF_INV_72\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_16\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[16]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_15_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[16]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_16_Z\, 
        CC => NET_CC_CONFIG152, P => NET_CC_CONFIG150, UB => 
        NET_CC_CONFIG151);
    
    \MemorySynchronizer_0/waitingtimercounter[13]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[13]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_53_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[13]\);
    
    \STAMP_0/un1_new_avail_0_sqmuxa_3\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/un1_new_avail_0_sqmuxa_1\, B => 
        \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_1\, Y => 
        \STAMP_0/un1_new_avail_0_sqmuxa_3_Z\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0_a2[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \MemorySynchronizer_0/un6_in_enable_i_0\, B
         => \MemorySynchronizer_0/MemorySyncState_Z[5]\, Y => 
        \MemorySynchronizer_0/N_1495\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_7\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[7]\, 
        B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_6_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_7_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_7_Z\, 
        CC => NET_CC_CONFIG648, P => NET_CC_CONFIG646, UB => 
        NET_CC_CONFIG647);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[15]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_76\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[15]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[15]\, 
        D => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[15]\);
    
    \MemorySynchronizer_0/MemorySyncState[1]\ : SLE
      port map(D => \MemorySynchronizer_0/MemorySyncState_ns[4]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, 
        EN => ENABLE_MEMORY_LED_c, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/MemorySyncState_Z[1]\);
    
    \STAMP_0/delay_counter_cry[0]_CC_0\ : CC_CONFIG
      port map(CI => ADLIB_GND0, CO => CI_TO_CO391, P(0) => 
        NET_CC_CONFIG393, P(1) => NET_CC_CONFIG396, P(2) => 
        NET_CC_CONFIG399, P(3) => NET_CC_CONFIG402, P(4) => 
        NET_CC_CONFIG405, P(5) => NET_CC_CONFIG408, P(6) => 
        NET_CC_CONFIG411, P(7) => NET_CC_CONFIG414, P(8) => 
        NET_CC_CONFIG417, P(9) => NET_CC_CONFIG420, P(10) => 
        NET_CC_CONFIG423, P(11) => NET_CC_CONFIG426, UB(0) => 
        NET_CC_CONFIG394, UB(1) => NET_CC_CONFIG397, UB(2) => 
        NET_CC_CONFIG400, UB(3) => NET_CC_CONFIG403, UB(4) => 
        NET_CC_CONFIG406, UB(5) => NET_CC_CONFIG409, UB(6) => 
        NET_CC_CONFIG412, UB(7) => NET_CC_CONFIG415, UB(8) => 
        NET_CC_CONFIG418, UB(9) => NET_CC_CONFIG421, UB(10) => 
        NET_CC_CONFIG424, UB(11) => NET_CC_CONFIG427, CC(0) => 
        NET_CC_CONFIG395, CC(1) => NET_CC_CONFIG398, CC(2) => 
        NET_CC_CONFIG401, CC(3) => NET_CC_CONFIG404, CC(4) => 
        NET_CC_CONFIG407, CC(5) => NET_CC_CONFIG410, CC(6) => 
        NET_CC_CONFIG413, CC(7) => NET_CC_CONFIG416, CC(8) => 
        NET_CC_CONFIG419, CC(9) => NET_CC_CONFIG422, CC(10) => 
        NET_CC_CONFIG425, CC(11) => NET_CC_CONFIG428);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a1\ : 
        CFG4
      generic map(INIT => x"2000")

      port map(A => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a1_0_Z\, 
        B => \sb_sb_0_STAMP_PADDR[5]\, C => 
        \MemorySynchronizer_0/N_271\, D => 
        \MemorySynchronizer_0/N_2564\, Y => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a1_Z\);
    
    \STAMP_0/dummy[0]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_40\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[0]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_10\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[10]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_9_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_10_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_10_Z\, CC
         => NET_CC_CONFIG755, P => NET_CC_CONFIG753, UB => 
        NET_CC_CONFIG754);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[3]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[3]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[3]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[3]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[11]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[11]\, B => 
        \sb_sb_0_STAMP_PWDATA[11]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[11]\);
    
    \STAMP_0/PRDATA[26]\ : SLE
      port map(D => \STAMP_0/N_676\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_41\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[26]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_66\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[10]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[10]\, B => 
        \sb_sb_0_STAMP_PWDATA[10]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[10]\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO_4[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[0]\, 
        B => \MemorySynchronizer_0/numberofnewavails_Z[1]\, Y => 
        \MemorySynchronizer_0/m3_e_0_0\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_20\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[20]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[20]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_19\, S => 
        \MemorySynchronizer_0/temp_1[20]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_20\, CC => 
        NET_CC_CONFIG259, P => NET_CC_CONFIG257, UB => 
        NET_CC_CONFIG258);
    
    \MemorySynchronizer_0/PREADY\ : SLE
      port map(D => \MemorySynchronizer_0/N_301\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => sb_sb_0_Memory_PREADY);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_166\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[29]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[29]\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/N_2323\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[29]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[29]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_RNIJ3231\ : 
        CFG4
      generic map(INIT => x"8ACF")

      port map(A => sb_sb_0_STAMP_PREADY, B => 
        sb_sb_0_Memory_PREADY, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/PREADY_0_iv_i\);
    
    \STAMP_0/measurement_temp[4]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[20]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_264\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net\);
    
    \STAMP_0/un45_async_state_cry_1\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \STAMP_0/config_Z[25]\, B => 
        \STAMP_0_data_frame[4]\, C => ADLIB_GND0, D => ADLIB_GND0, 
        FCI => \STAMP_0/un45_async_state_cry_0_Z\, S => OPEN, Y
         => OPEN, FCO => \STAMP_0/un45_async_state_cry_1_Z\, CC
         => NET_CC_CONFIG519, P => NET_CC_CONFIG517, UB => 
        NET_CC_CONFIG518);
    
    \STAMP_0/component_state[2]\ : SLE
      port map(D => \STAMP_0/component_state_ns[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/component_state_Z[2]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_37_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[23]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_37\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO_1[5]\ : CFG4
      generic map(INIT => x"0A08")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[5]\, B
         => \MemorySynchronizer_0/g2_0_0\, C => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, D => 
        \MemorySynchronizer_0/g3\, Y => \MemorySynchronizer_0/g2\);
    
    \STAMP_0/un45_async_state_cry_5_FCINST1\ : FCEND_BUFF_CC
      port map(FCI => \STAMP_0/un45_async_state_cry_5_FCNET1\, CO
         => \STAMP_0/un45_async_state_cry_5_Z\, CC => 
        NET_CC_CONFIG534, P => NET_CC_CONFIG532, UB => 
        NET_CC_CONFIG533);
    
    \STAMP_0/delay_counter_s[27]\ : ARI1_CC
      generic map(INIT => x"45500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[27]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[26]\, S
         => \STAMP_0/delay_counter_s_Z[27]\, Y => OPEN, FCO => 
        OPEN, CC => NET_CC_CONFIG476, P => NET_CC_CONFIG474, UB
         => NET_CC_CONFIG475);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[10]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[10]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[9]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[10]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[10]\, CC
         => NET_CC_CONFIG36, P => NET_CC_CONFIG34, UB => 
        NET_CC_CONFIG35);
    
    \STAMP_0/un1_spi_rx_data_1[15]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[47]\, B => 
        \STAMP_0/dummy_Z[15]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_632\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_287\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[24]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_24_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[8]\);
    
    \STAMP_0/PRDATA[4]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[4]\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO_2[5]\ : CFG3
      generic map(INIT => x"02")

      port map(A => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, B
         => STAMP_0_new_avail, C => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[15]\, Y
         => \MemorySynchronizer_0/SynchStatusReg_RNO_2_Z[5]\);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_30_FCINST1\ : 
        FCEND_BUFF_CC
      port map(FCI => 
        \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_30_FCNET1\, 
        CO => \MemorySynchronizer_0/temp_1_cry_30\, CC => 
        NET_CC_CONFIG292, P => NET_CC_CONFIG290, UB => 
        NET_CC_CONFIG291);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_5\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_6\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_4_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[6]\, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_5_Z\, 
        CC => NET_CC_CONFIG1038, P => NET_CC_CONFIG1036, UB => 
        NET_CC_CONFIG1037);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[1]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[1]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1[31]\, Y => 
        \MemorySynchronizer_0/N_1090\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[0]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[0]\, 
        B => \MemorySynchronizer_0/un1_MemorySyncState_11_i\, C
         => ENABLE_MEMORY_LED_c, D => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[32]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[21]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[21]\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0[2]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => STAMP_0_new_avail, C => 
        \MemorySynchronizer_0/N_1495\, D => 
        \MemorySynchronizer_0/N_140_2\, Y => 
        \MemorySynchronizer_0/MemorySyncState_ns[2]\);
    
    \MemorySynchronizer_0/ConfigReg[18]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[18]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_44\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[16]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_44_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[6]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[6]\);
    
    \MemorySynchronizer_0/SynchStatusReg[23]\ : SLE
      port map(D => \MemorySynchronizer_0/N_2032_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[23]\);
    
    \MemorySynchronizer_0/end_one_counter_RNO[0]\ : CFG3
      generic map(INIT => x"C1")

      port map(A => \MemorySynchronizer_0/end_one_counter_Z[1]\, 
        B => \MemorySynchronizer_0/N_2337\, C => 
        \MemorySynchronizer_0/end_one_counter_Z[0]\, Y => 
        \MemorySynchronizer_0/N_207_i\);
    
    \MemorySynchronizer_0/SynchStatusReg2_RNO[11]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \MemorySynchronizer_0/temp_1_cry_0_Y\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[11]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[11]\);
    
    \STAMP_0/un1_spi_rx_data[14]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_664\, C => \STAMP_0/spi_rx_data[14]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[14]\);
    
    \STAMP_0/status_async_cycles_3_sqmuxa_0_a3\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_1\, 
        B => \STAMP_0/async_state_Z[1]\, C => 
        \STAMP_0/un1_async_prescaler_count\, Y => 
        \STAMP_0/status_async_cycles_3_sqmuxa\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_30\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un104_in_enable_30\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[30]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_29_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_30_Z\, CC => 
        NET_CC_CONFIG913, P => NET_CC_CONFIG911, UB => 
        NET_CC_CONFIG912);
    
    \MemorySynchronizer_0/resynctimercounter[23]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1099\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[23]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[16]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_16\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[16]\, 
        C => \MemorySynchronizer_0/N_1517\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[16]\);
    
    \MemorySynchronizer_0/resettimercounter[26]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_28_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[26]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_34\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg2_RNO[9]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[3]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[9]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[9]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[8]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[2]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[8]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[8]\);
    
    AFLSDF_INV_38 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_38\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[17]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[17]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1074\, Y => 
        \MemorySynchronizer_0/N_1105\);
    
    \STAMP_0/spi/count_cry[24]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[24]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[23]\, S => 
        \STAMP_0/spi/count_s[24]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[24]\, CC => NET_CC_CONFIG997, P
         => NET_CC_CONFIG995, UB => NET_CC_CONFIG996);
    
    \STAMP_0/PRDATA_RNO[30]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => \STAMP_0/N_220\, B => \STAMP_0/N_218\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_5\, D => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_119_i\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[23]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[23]\, B => 
        \sb_sb_0_STAMP_PWDATA[23]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[23]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_46\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[7]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_ResetTimerValueReg_46_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_236\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46]\, 
        IPC => OPEN);
    
    AFLSDF_INV_49 : INV_BA
      port map(A => NN_1, Y => \AFLSDF_INV_49\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_CC_1\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO100, CO => CI_TO_CO101, P(0) => 
        NET_CC_CONFIG135, P(1) => NET_CC_CONFIG138, P(2) => 
        NET_CC_CONFIG141, P(3) => NET_CC_CONFIG144, P(4) => 
        NET_CC_CONFIG147, P(5) => NET_CC_CONFIG150, P(6) => 
        NET_CC_CONFIG153, P(7) => NET_CC_CONFIG156, P(8) => 
        NET_CC_CONFIG159, P(9) => NET_CC_CONFIG162, P(10) => 
        NET_CC_CONFIG165, P(11) => NET_CC_CONFIG168, UB(0) => 
        NET_CC_CONFIG136, UB(1) => NET_CC_CONFIG139, UB(2) => 
        NET_CC_CONFIG142, UB(3) => NET_CC_CONFIG145, UB(4) => 
        NET_CC_CONFIG148, UB(5) => NET_CC_CONFIG151, UB(6) => 
        NET_CC_CONFIG154, UB(7) => NET_CC_CONFIG157, UB(8) => 
        NET_CC_CONFIG160, UB(9) => NET_CC_CONFIG163, UB(10) => 
        NET_CC_CONFIG166, UB(11) => NET_CC_CONFIG169, CC(0) => 
        NET_CC_CONFIG137, CC(1) => NET_CC_CONFIG140, CC(2) => 
        NET_CC_CONFIG143, CC(3) => NET_CC_CONFIG146, CC(4) => 
        NET_CC_CONFIG149, CC(5) => NET_CC_CONFIG152, CC(6) => 
        NET_CC_CONFIG155, CC(7) => NET_CC_CONFIG158, CC(8) => 
        NET_CC_CONFIG161, CC(9) => NET_CC_CONFIG164, CC(10) => 
        NET_CC_CONFIG167, CC(11) => NET_CC_CONFIG170);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_104\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[4]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg[25]\ : SLE
      port map(D => \MemorySynchronizer_0/N_2033_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[25]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_188\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/status_async_cycles_lm_0[5]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/status_async_cycles_3_sqmuxa\, B => 
        \STAMP_0/status_async_cycles_s_Z[5]\, C => 
        \STAMP_0/status_async_cycles_1_sqmuxa_Z\, Y => 
        \STAMP_0/status_async_cycles_lm[5]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[17]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[17]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[16]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[17]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[17]\, CC
         => NET_CC_CONFIG57, P => NET_CC_CONFIG55, UB => 
        NET_CC_CONFIG56);
    
    \MemorySynchronizer_0/resettimercounter[28]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_19_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[28]\);
    
    AFLSDF_INV_47 : INV_BA
      port map(A => \MemorySynchronizer_0/N_1981_i\, Y => 
        \AFLSDF_INV_47\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_23\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_24\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_22_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[24]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_23_Z\, CC
         => NET_CC_CONFIG1092, P => NET_CC_CONFIG1090, UB => 
        NET_CC_CONFIG1091);
    
    \MemorySynchronizer_0/un104_in_enable_cry_14\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[14]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[14]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_13_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_14_Z\, CC => 
        NET_CC_CONFIG865, P => NET_CC_CONFIG863, UB => 
        NET_CC_CONFIG864);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[5]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[5]\, 
        B => \sb_sb_0_STAMP_PWDATA[5]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[5]\);
    
    \STAMP_0/un1_PREADY_0_sqmuxa_3_0_RNO\ : CFG2
      generic map(INIT => x"4")

      port map(A => sb_sb_0_STAMP_PENABLE, B => 
        \STAMP_0/component_state_Z[2]\, Y => \STAMP_0/N_162_i\);
    
    \STAMP_0/un1_spi_rx_data_2[9]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_592\, B => \STAMP_0/N_626\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_659\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[28]\ : SLE
      port map(D => \STAMP_0_data_frame[60]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[28]\);
    
    \MemorySynchronizer_0/resettimercounter[21]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_12_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[21]\);
    
    \STAMP_0/config[20]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[20]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[16]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[16]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_9[28]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_2569\, C => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_2577\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_232\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[1]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[1]\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_21_Z\, B => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_20_Z\, C => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_27_Z\, D => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_28_Z\, Y => 
        \MemorySynchronizer_0/un6_in_enable_i_0\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_19\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/N_1078\, B => 
        \MemorySynchronizer_0/N_1077\, C => 
        \MemorySynchronizer_0/N_1062\, D => 
        \MemorySynchronizer_0/N_1061\, Y => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_19_Z\);
    
    \STAMP_0/spi/tx_buffer_RNO[5]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[5]\, B => 
        \STAMP_0/spi/tx_buffer_Z[4]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_132\);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_16\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[7]\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[6]\, C => 
        \MemorySynchronizer_0/waitingtimercounter_Z[4]\, D => 
        \MemorySynchronizer_0/waitingtimercounter_Z[1]\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_16_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1[4]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_0_Z[4]\, 
        B => \MemorySynchronizer_0/N_2510\, C => 
        \MemorySynchronizer_0/SynchStatusReg_Z[6]\, D => 
        \MemorySynchronizer_0/N_2606\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168[4]\);
    
    \MemorySynchronizer_0/ConfigReg[24]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[24]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_16\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[16]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_15_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_16_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_16_Z\, 
        CC => NET_CC_CONFIG675, P => NET_CC_CONFIG673, UB => 
        NET_CC_CONFIG674);
    
    \STAMP_0/spi/rx_data[6]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[6]\);
    
    \MemorySynchronizer_0/un1_nreset_16_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_43_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_16_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_16_rs_Z\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_26\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[26]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_25_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_26_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_26_Z\, CC
         => NET_CC_CONFIG803, P => NET_CC_CONFIG801, UB => 
        NET_CC_CONFIG802);
    
    \STAMP_0/spi_dms1_cs_0_sqmuxa_3_0_a3\ : CFG3
      generic map(INIT => x"80")

      port map(A => \STAMP_0/drdy_flank_detected_dms1_Z\, B => 
        \STAMP_0/config_Z[30]\, C => \STAMP_0/N_333\, Y => 
        \STAMP_0/spi_dms1_cs_0_sqmuxa_3\);
    
    \MemorySynchronizer_0/TimeStampReg[9]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[9]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[9]\);
    
    \STAMP_0/un1_spi_rx_data[10]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_660\, C => \STAMP_0/spi_rx_data[10]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[10]\);
    
    \STAMP_0/spi/count[18]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[18]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_260\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[9]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_9_S\, 
        Y => \MemorySynchronizer_0/N_1533\);
    
    \MemorySynchronizer_0/SynchStatusReg2[23]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[23]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[25]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[25]\, B => 
        \sb_sb_0_Memory_PRDATA[25]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[25]\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0_a3_0[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/MemorySyncState_Z[2]\, Y => 
        \MemorySynchronizer_0/N_1482\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[10]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[10]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[10]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[22]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[10]\);
    
    \STAMP_0/spi/rx_buffer[8]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[8]\);
    
    \STAMP_0/request_resync_0_sqmuxa_0_a3\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/component_state_Z[5]\, B => 
        \STAMP_0/config_Z[31]\, Y => 
        \STAMP_0/request_resync_0_sqmuxa\);
    
    \stamp0_ready_dms1_ibuf/U0/U_IOIN\ : IOIN_IB
      port map(YIN => \stamp0_ready_dms1_ibuf/U0/YIN\, E => 
        ADLIB_GND0, Y => stamp0_ready_dms1_c);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[6]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[6]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[6]\, C => 
        \MemorySynchronizer_0/N_2596\, D => 
        \MemorySynchronizer_0/N_2595\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[6]\);
    
    \MemorySynchronizer_0/TimeStampReg[21]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[21]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[21]\);
    
    \MemorySynchronizer_0/waitingtimercounter[25]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[25]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_26_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[25]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[4]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_4\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[4]\, 
        C => \MemorySynchronizer_0/N_1549\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[4]\);
    
    \STAMP_0/spi/count_cry[8]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[8]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[7]\, S => 
        \STAMP_0/spi/count_s[8]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[8]\, CC => NET_CC_CONFIG949, P
         => NET_CC_CONFIG947, UB => NET_CC_CONFIG948);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_1[11]\ : CFG4
      generic map(INIT => x"00E0")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[13]\, 
        B => \STAMP_0_data_frame[9]\, C => 
        \MemorySynchronizer_0/MemorySyncState_Z[5]\, D => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_1_Z[11]\);
    
    \STAMP_0/async_prescaler_count[5]\ : SLE
      port map(D => \STAMP_0/un5_async_prescaler_count_cry_5_S\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[5]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[11]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_11\);
    
    \STAMP_0/spi/tx_buffer_RNO[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[8]\, B => 
        \STAMP_0/spi/tx_buffer_Z[7]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_127\);
    
    \STAMP_0/async_prescaler_count[6]\ : SLE
      port map(D => \STAMP_0/async_prescaler_count_5_Z[6]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[6]\);
    
    \STAMP_0/spi/count[5]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[5]\);
    
    \STAMP_0/spi/count[27]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[27]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[16]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[16]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[15]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[16]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[16]\, CC
         => NET_CC_CONFIG54, P => NET_CC_CONFIG52, UB => 
        NET_CC_CONFIG53);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_9\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[9]\, 
        B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_8_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_9_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_9_Z\, 
        CC => NET_CC_CONFIG654, P => NET_CC_CONFIG652, UB => 
        NET_CC_CONFIG653);
    
    \MemorySynchronizer_0/SynchStatusReg2[17]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[17]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[17]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_10\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[10]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_9_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[10]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_10_Z\, 
        CC => NET_CC_CONFIG134, P => NET_CC_CONFIG132, UB => 
        NET_CC_CONFIG133);
    
    \MemorySynchronizer_0/un1_nreset_56_0_a3_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[10]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_56_i\);
    
    \STAMP_0/un1_spi_rx_data_2[31]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_614\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, C => \STAMP_0/N_648\, Y
         => \STAMP_0/N_681\);
    
    \STAMP_0/un1_spi_rx_data_2[28]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_611\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, C => \STAMP_0/N_645\, Y
         => \STAMP_0/N_678\);
    
    AFLSDF_INV_23 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_23\);
    
    \LED_RECORDING_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \LED_RECORDING_obuf/U0/DOUT1\, Y => 
        \LED_RECORDING_obuf/U0/DOUT\);
    
    AFLSDF_INV_83 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_83\);
    
    \MOSI_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \MOSI_obuf/U0/EOUT1\, Y => 
        \MOSI_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_0_CC_1\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO721, CO => CI_TO_CO722, P(0) => 
        NET_CC_CONFIG759, P(1) => NET_CC_CONFIG762, P(2) => 
        NET_CC_CONFIG765, P(3) => NET_CC_CONFIG768, P(4) => 
        NET_CC_CONFIG771, P(5) => NET_CC_CONFIG774, P(6) => 
        NET_CC_CONFIG777, P(7) => NET_CC_CONFIG780, P(8) => 
        NET_CC_CONFIG783, P(9) => NET_CC_CONFIG786, P(10) => 
        NET_CC_CONFIG789, P(11) => NET_CC_CONFIG792, UB(0) => 
        NET_CC_CONFIG760, UB(1) => NET_CC_CONFIG763, UB(2) => 
        NET_CC_CONFIG766, UB(3) => NET_CC_CONFIG769, UB(4) => 
        NET_CC_CONFIG772, UB(5) => NET_CC_CONFIG775, UB(6) => 
        NET_CC_CONFIG778, UB(7) => NET_CC_CONFIG781, UB(8) => 
        NET_CC_CONFIG784, UB(9) => NET_CC_CONFIG787, UB(10) => 
        NET_CC_CONFIG790, UB(11) => NET_CC_CONFIG793, CC(0) => 
        NET_CC_CONFIG761, CC(1) => NET_CC_CONFIG764, CC(2) => 
        NET_CC_CONFIG767, CC(3) => NET_CC_CONFIG770, CC(4) => 
        NET_CC_CONFIG773, CC(5) => NET_CC_CONFIG776, CC(6) => 
        NET_CC_CONFIG779, CC(7) => NET_CC_CONFIG782, CC(8) => 
        NET_CC_CONFIG785, CC(9) => NET_CC_CONFIG788, CC(10) => 
        NET_CC_CONFIG791, CC(11) => NET_CC_CONFIG794);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_51\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[7]\, 
        B => \MemorySynchronizer_0/un104_in_enable_6\, C => 
        \MemorySynchronizer_0/un104_in_enable_7\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[6]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[2]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[3]\, CC
         => NET_CC_CONFIG547, P => NET_CC_CONFIG545, UB => 
        NET_CC_CONFIG546);
    
    \LED_RECORDING_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => LED_RECORDING, D => 
        \LED_RECORDING_obuf/U0/DOUT\, E => 
        \LED_RECORDING_obuf/U0/EOUT\);
    
    \STAMP_0/delay_counter_cry[25]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[25]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[24]\, S
         => \STAMP_0/delay_counter_s[25]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[25]\, CC => NET_CC_CONFIG470, 
        P => NET_CC_CONFIG468, UB => NET_CC_CONFIG469);
    
    \STAMP_0/config[5]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[5]\);
    
    \STAMP_0/delay_counter_cry[4]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[4]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/delay_counter_cry_Z[3]\, S => 
        \STAMP_0/delay_counter_s[4]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[4]\, CC => NET_CC_CONFIG407, 
        P => NET_CC_CONFIG405, UB => NET_CC_CONFIG406);
    
    \STAMP_0/spi_tx_data_RNO[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[3]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_295_i\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_20\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_16_S\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_17_S\, 
        C => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_18_S\, D
         => \MemorySynchronizer_0/un5_resettimercounter_cry_19_S\, 
        Y => \MemorySynchronizer_0/un6_in_enable_0_a3_20_Z\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[11]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[11]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[21]\, Y
         => \MemorySynchronizer_0/N_1080\);
    
    \STAMP_0/measurement_dms2[14]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[46]\);
    
    AFLSDF_INV_14 : INV_BA
      port map(A => \sb_sb_0/CCC_0/GL1_net\, Y => \AFLSDF_INV_14\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_40_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_42\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_40_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_53\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14]\, 
        IPC => OPEN);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB0\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB0_rgbr_net_1\);
    
    \STAMP_0/spi/rx_buffer[15]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[15]\);
    
    \resetn_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \resetn_obuf/U0/EOUT1\, Y => 
        \resetn_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_0\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[0]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => ADLIB_GND0, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_0_Z\, CC
         => NET_CC_CONFIG297, P => NET_CC_CONFIG295, UB => 
        NET_CC_CONFIG296);
    
    \debug_led_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => ADLIB_GND0, E => ADLIB_VCC1, DOUT => 
        \debug_led_obuf/U0/DOUT1\, EOUT => 
        \debug_led_obuf/U0/EOUT1\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[10]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[10]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[10]\);
    
    \STAMP_0/dummy[1]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_43\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[1]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_127\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9]\, 
        IPC => OPEN);
    
    \STAMP_0/measurement_dms2[11]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[43]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_25\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[25]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_24_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_25_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_25_Z\, CC
         => NET_CC_CONFIG800, P => NET_CC_CONFIG798, UB => 
        NET_CC_CONFIG799);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_21\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[18]\, B => 
        \MemorySynchronizer_0/un120_in_enable_i_A[19]\, C => 
        \MemorySynchronizer_0/un120_in_enable_i_A[20]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[21]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_21_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_73\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/TimeStampReg[11]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[11]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[11]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[12]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_12_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_72\);
    
    AFLSDF_INV_26 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_26\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_10\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[10]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[10]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_9_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_10_Z\, CC => 
        NET_CC_CONFIG853, P => NET_CC_CONFIG851, UB => 
        NET_CC_CONFIG852);
    
    \STAMP_0/spi/count_lm_0[2]\ : CFG4
      generic map(INIT => x"D8CC")

      port map(A => \STAMP_0/spi/un7_count_NE_i\, B => 
        \STAMP_0/spi/count_0_sqmuxa\, C => 
        \STAMP_0/spi/count_s[2]\, D => \STAMP_0/spi/state_Z[0]\, 
        Y => \STAMP_0/spi/count_lm[2]\);
    
    \MemorySynchronizer_0/SynchStatusReg[30]\ : SLE
      port map(D => \MemorySynchronizer_0/N_2015_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[30]\);
    
    \STAMP_0/spi/busy_RNIS7HJ\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/component_state_Z[0]\, B => 
        \STAMP_0/spi_busy\, Y => \STAMP_0/N_353\);
    
    \STAMP_0/measurement_dms2[5]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[37]\);
    
    AFLSDF_INV_86 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_86\);
    
    \MemorySynchronizer_0/un1_nreset_13\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[20]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_13_i\);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.un151_in_enablelto30_16\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/temp_1[17]\, B => 
        \MemorySynchronizer_0/temp_1[18]\, C => 
        \MemorySynchronizer_0/temp_1[19]\, D => 
        \MemorySynchronizer_0/temp_1[20]\, Y => 
        \MemorySynchronizer_0/un151_in_enablelto30_16\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[16]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[16]\, B => 
        \sb_sb_0_STAMP_PWDATA[16]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[16]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_22\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[22]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_21_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_22_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_22_Z\, 
        CC => NET_CC_CONFIG693, P => NET_CC_CONFIG691, UB => 
        NET_CC_CONFIG692);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4[8]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \MemorySynchronizer_0/un104_in_enable_8\, B
         => \MemorySynchronizer_0/SynchStatusReg2_Z[8]\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2594\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[8]\);
    
    \STAMP_0/async_prescaler_count[7]\ : SLE
      port map(D => \STAMP_0/async_prescaler_count_5_Z[7]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[7]\);
    
    \MemorySynchronizer_0/resettimercounter[12]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_41_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[12]\);
    
    \MemorySynchronizer_0/un1_nreset_42_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_50\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_42_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_42_rs_Z\);
    
    \MemorySynchronizer_0/un1_nreset_36_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_43\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_36_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_36_rs_Z\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[7]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_7\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_34_RNO_0[20]\ : 
        CFG3
      generic map(INIT => x"7F")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[2]\, 
        B => \MemorySynchronizer_0/numberofnewavails_Z[1]\, C => 
        \MemorySynchronizer_0/numberofnewavails_Z[0]\, Y => 
        \MemorySynchronizer_0/g0_0_1\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[4]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[4]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1087\, Y => 
        \MemorySynchronizer_0/N_1118\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[17]\ : SLE
      port map(D => \STAMP_0_data_frame[49]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[17]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_o2[4]\ : CFG4
      generic map(INIT => x"4F0F")

      port map(A => \MemorySynchronizer_0/N_2313\, B => 
        \MemorySynchronizer_0/N_140_1_i\, C => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_o2_1_0[4]\, 
        D => \MemorySynchronizer_0/N_140_2\, Y => 
        \MemorySynchronizer_0/N_2326\);
    
    \MemorySynchronizer_0/resettimercounter_RNI7Q6V[21]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_1980_i_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[21]\, C => 
        \MemorySynchronizer_0/un1_nreset_12_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[21]\);
    
    \STAMP_0/spi/count_cry[26]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[26]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[25]\, S => 
        \STAMP_0/spi/count_s[26]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[26]\, CC => NET_CC_CONFIG1003, P
         => NET_CC_CONFIG1001, UB => NET_CC_CONFIG1002);
    
    \STAMP_0/apb_spi_finished_1_sqmuxa_0_a3\ : CFG3
      generic map(INIT => x"80")

      port map(A => \STAMP_0/spi_request_for_Z[1]\, B => 
        \STAMP_0/spi_request_for_Z[0]\, C => 
        \STAMP_0/apb_spi_finished_0_sqmuxa_1\, Y => 
        \STAMP_0/apb_spi_finished_1_sqmuxa\);
    
    \MMUART_0_TXD_M2F_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \MMUART_0_TXD_M2F_obuf/U0/EOUT1\, Y => 
        \MMUART_0_TXD_M2F_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/un1_nreset_27_rs_RNI7I3N\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_55_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[27]\, C => 
        \MemorySynchronizer_0/un1_nreset_27_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[27]\);
    
    \STAMP_0/spi/clk_toggles[2]\ : SLE
      port map(D => \STAMP_0/spi/clk_toggles_lm[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB14_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_37_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/clk_toggles_Z[2]\);
    
    \MemorySynchronizer_0/resynctimercounter[1]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1121\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[1]\);
    
    \STAMP_0/delay_counter_cry[5]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[5]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/delay_counter_cry_Z[4]\, S => 
        \STAMP_0/delay_counter_s[5]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[5]\, CC => NET_CC_CONFIG410, 
        P => NET_CC_CONFIG408, UB => NET_CC_CONFIG409);
    
    \MemorySynchronizer_0/ResetTimerValueReg[9]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[9]\);
    
    \STAMP_0/async_prescaler_count_5[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/un1_async_prescaler_count\, B => 
        \STAMP_0/un5_async_prescaler_count_cry_7_S\, Y => 
        \STAMP_0/async_prescaler_count_5_Z[7]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_FCINST1\ : 
        FCEND_BUFF_CC
      port map(FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_FCNET1\, 
        CO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_Z\, 
        CC => NET_CC_CONFIG1113, P => NET_CC_CONFIG1111, UB => 
        NET_CC_CONFIG1112);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[16]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[16]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[16]\, Y
         => \MemorySynchronizer_0/N_1075\);
    
    \STAMP_0/delay_counter_lm_0[27]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s_Z[27]\, Y => 
        \STAMP_0/delay_counter_lm[27]\);
    
    \STAMP_0/delay_counter_cry[6]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[6]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/delay_counter_cry_Z[5]\, S => 
        \STAMP_0/delay_counter_s[6]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[6]\, CC => NET_CC_CONFIG413, 
        P => NET_CC_CONFIG411, UB => NET_CC_CONFIG412);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[19]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[19]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[19]\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[19]\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[19]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_19\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[19]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_18_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[19]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_19_Z\, 
        CC => NET_CC_CONFIG161, P => NET_CC_CONFIG159, UB => 
        NET_CC_CONFIG160);
    
    \STAMP_0/spi/assert_data_5_iv_0_0\ : CFG4
      generic map(INIT => x"52A2")

      port map(A => \STAMP_0/spi/assert_data_Z\, B => 
        \STAMP_0/enable\, C => \STAMP_0/spi/state_Z[0]\, D => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/assert_data_5\);
    
    \STAMP_0/spi/un7_count_NE_27\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \STAMP_0/spi/count_Z[26]\, B => 
        \STAMP_0/spi/count_Z[27]\, C => 
        \STAMP_0/spi/un7_count_NE_23_Z\, D => 
        \STAMP_0/spi/un7_count_NE_13_Z\, Y => 
        \STAMP_0/spi/un7_count_NE_27_Z\);
    
    \STAMP_0/delay_counter_cry[0]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[0]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => ADLIB_GND0, S
         => OPEN, Y => \STAMP_0/delay_counter_cry_Y[0]\, FCO => 
        \STAMP_0/delay_counter_cry_Z[0]\, CC => NET_CC_CONFIG395, 
        P => NET_CC_CONFIG393, UB => NET_CC_CONFIG394);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[7]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[7]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[13]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_13_S\, 
        Y => \MemorySynchronizer_0/N_1525\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[3]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[3]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[29]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[3]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[29]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[29]\);
    
    \STAMP_0/config[25]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[25]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_52_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[14]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_52\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[10]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_10_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[22]\);
    
    \STAMP_0/request_resync\ : SLE
      port map(D => \STAMP_0/request_resync_1_sqmuxa_1_Z\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN
         => \STAMP_0/N_152\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[9]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_28[20]\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_2_Z[20]\, 
        B => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_14_Z[20]\, 
        C => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_25_Z[20]\, 
        D => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_21_Z[20]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_28_Z[20]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_231\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41]\, 
        IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data_0[26]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame[26]\, B => 
        \STAMP_0/config_Z[26]\, C => \sb_sb_0_STAMP_PADDR[8]\, Y
         => \STAMP_0/N_609\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[6]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[6]\, B => 
        \sb_sb_0_Memory_PRDATA[6]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6]\);
    
    \MemorySynchronizer_0/dataReadyReset_RNO\ : CFG4
      generic map(INIT => x"030A")

      port map(A => MemorySynchronizer_0_dataReadyReset, B => 
        \MemorySynchronizer_0/end_one_counter_Z[1]\, C => 
        \MemorySynchronizer_0/MemorySyncState_Z[5]\, D => 
        \MemorySynchronizer_0/MemorySyncState_Z[1]\, Y => 
        \MemorySynchronizer_0/N_2068_i\);
    
    \STAMP_0/delay_counter[27]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[27]\);
    
    \MemorySynchronizer_0/TimeStampReg[22]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[22]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[22]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[29]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[29]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_29\);
    
    \MemorySynchronizer_0/un94_in_enable_18\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[26]\, B => 
        \MemorySynchronizer_0/resettimercounter_Z[25]\, C => 
        \MemorySynchronizer_0/resettimercounter_Z[24]\, D => 
        \MemorySynchronizer_0/resettimercounter_Z[23]\, Y => 
        \MemorySynchronizer_0/un94_in_enable_18_Z\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_42_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_44\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_42_set_Z\);
    
    \MemorySynchronizer_0/resettimercounter[7]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[7]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_48_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[7]\);
    
    \STAMP_0/drdy_flank_detected_temp\ : SLE
      port map(D => \STAMP_0/stamp0_ready_temp_c_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_2_i_Z\, ALn
         => \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/drdy_flank_detected_temp_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[28]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[28]\, B => 
        \sb_sb_0_STAMP_PWDATA[28]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[28]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[22]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_22_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[10]\);
    
    \MemorySynchronizer_0/N_2532_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_45\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_2532_set_Z\);
    
    \STAMP_0/async_prescaler_count[2]\ : SLE
      port map(D => \STAMP_0/async_prescaler_count_5_Z[2]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[2]\);
    
    \MemorySynchronizer_0/N_1979_i_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_46\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_1979_i_set_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[30]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[30]\, B => 
        \MemorySynchronizer_0/un104_in_enable_30\, C => 
        \MemorySynchronizer_0/N_2574\, D => 
        \MemorySynchronizer_0/N_2577\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[30]\);
    
    \STAMP_0/un1_component_state_14_i_a3_0_2\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/N_337\, B => 
        \STAMP_0/spi_request_for_Z[1]\, C => \STAMP_0/N_331\, Y
         => \STAMP_0/N_248_2\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[1]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[1]\);
    
    \STAMP_0/measurement_dms1[12]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[60]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[3]\ : SLE
      port map(D => \STAMP_0_data_frame[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[3]\);
    
    \MemorySynchronizer_0/N_2533_set_RNI9RF41\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_2533_set_Z\, B => 
        \MemorySynchronizer_0/waitingtimercounterrs[9]\, C => 
        \MemorySynchronizer_0/un1_nreset_57_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[9]\);
    
    \MemorySynchronizer_0/SynchStatusReg[31]\ : SLE
      port map(D => \MemorySynchronizer_0/N_2016_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[31]\);
    
    \STAMP_0/un5_async_prescaler_count_s_1_391\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[0]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => ADLIB_VCC1, S => OPEN, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_s_1_391_FCO\, 
        CC => NET_CC_CONFIG480, P => NET_CC_CONFIG478, UB => 
        NET_CC_CONFIG479);
    
    \ENABLE_MEMORY_LED_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => ENABLE_MEMORY_LED_c, E => ADLIB_VCC1, DOUT
         => \ENABLE_MEMORY_LED_obuf/U0/DOUT1\, EOUT => 
        \ENABLE_MEMORY_LED_obuf/U0/EOUT1\);
    
    \STAMP_0/un1_spi_rx_data_0[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[3]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[3]\, Y
         => \STAMP_0/N_586\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_157\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/measurement_dms1[3]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[51]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_35_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[18]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_35\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[8]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[8]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1083\, Y => 
        \MemorySynchronizer_0/N_1114\);
    
    \MemorySynchronizer_0/waitingtimercounter[24]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[24]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_42_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[24]\);
    
    \MemorySynchronizer_0/N_1981_i_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_47\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_1981_i_set_Z\);
    
    \STAMP_0/spi/count_lm_0[20]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[20]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[20]\);
    
    \STAMP_0/un1_spi_rx_data[12]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_662\, C => \STAMP_0/spi_rx_data[12]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[12]\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_13\ : CFG2
      generic map(INIT => x"1")

      port map(A => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_27_S\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_26_S\, 
        Y => \MemorySynchronizer_0/un6_in_enable_0_a3_13_Z\);
    
    \STAMP_0/spi/clk_toggles_lm_0[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/spi/ss_n_buffer_1_sqmuxa\, B => 
        \STAMP_0/spi/clk_toggles_s[2]\, Y => 
        \STAMP_0/spi/clk_toggles_lm[2]\);
    
    \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_2_i\ : CFG3
      generic map(INIT => x"FD")

      port map(A => stamp0_ready_dms2_c, B => 
        \STAMP_0/request_resync_0_sqmuxa\, C => 
        \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_1\, Y => 
        \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_2_i_Z\);
    
    \STAMP_0/delay_counter[3]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[3]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_18\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[18]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_17_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_18_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_18_Z\, 
        CC => NET_CC_CONFIG681, P => NET_CC_CONFIG679, UB => 
        NET_CC_CONFIG680);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_52_i_i_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[1]\, B => NN_1, 
        Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_52_i_i_a2_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_34[20]\ : 
        CFG4
      generic map(INIT => x"0A0E")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[22]\, 
        B => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_31_Z[20]\, 
        C => \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, D
         => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_34_1[20]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_34_Z[20]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[25]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[25]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[7]\, Y => 
        \MemorySynchronizer_0/N_1066\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_33_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_48\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_33_set_Z\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_43_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[29]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_43\);
    
    \STAMP_0/spi/count_lm_0[5]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[5]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[5]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_267\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un104_in_enable_cry_17\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[17]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[17]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_16_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_17_Z\, CC => 
        NET_CC_CONFIG874, P => NET_CC_CONFIG872, UB => 
        NET_CC_CONFIG873);
    
    \STAMP_0/apb_is_atomic_0_sqmuxa_0_a3\ : CFG2
      generic map(INIT => x"8")

      port map(A => debug_led_net_0, B => 
        \STAMP_0/apb_spi_finished_0_sqmuxa\, Y => 
        \STAMP_0/apb_is_atomic_0_sqmuxa\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[11]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[11]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1080\, Y => 
        \MemorySynchronizer_0/N_1111\);
    
    AFLSDF_INV_59 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_39\, Y => 
        \AFLSDF_INV_59\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_17\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[2]\, 
        B => \MemorySynchronizer_0/un120_in_enable_i_A[5]\, C => 
        \MemorySynchronizer_0/un120_in_enable_i_A[4]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[3]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_17_Z\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_1\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[1]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[1]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_0\, S => 
        \MemorySynchronizer_0/temp_1[1]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_1\, CC => 
        NET_CC_CONFIG202, P => NET_CC_CONFIG200, UB => 
        NET_CC_CONFIG201);
    
    \STAMP_0/config_RNO[31]\ : CFG4
      generic map(INIT => x"E222")

      port map(A => \STAMP_0/component_state_Z[5]\, B => 
        \STAMP_0/component_state_Z[3]\, C => \STAMP_0/un76_paddr\, 
        D => sb_sb_0_STAMP_PWRITE, Y => 
        \STAMP_0/un1_component_state_6_i\);
    
    \STAMP_0/delay_counter_RNI20MA[16]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \STAMP_0/delay_counter_Z[19]\, B => 
        \STAMP_0/delay_counter_Z[18]\, C => 
        \STAMP_0/delay_counter_Z[17]\, D => 
        \STAMP_0/delay_counter_Z[16]\, Y => 
        \STAMP_0/N_517_i_0_a2_14\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[25]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[25]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[25]\, D
         => \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[25]\);
    
    \MemorySynchronizer_0/TimeStampReg[12]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[12]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[12]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[29]\ : SLE
      port map(D => \STAMP_0_data_frame[61]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[29]\);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_20\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[29]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[27]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[26]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[25]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_20_Z\);
    
    \STAMP_0/spi/count_lm_0[28]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[28]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[28]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_27[20]\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_18_Z[20]\, 
        B => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_17_Z[20]\, 
        C => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_16_Z[20]\, 
        D => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_15_Z[20]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_27_Z[20]\);
    
    AFLSDF_INV_57 : INV_BA
      port map(A => \MemorySynchronizer_0/N_21_i\, Y => 
        \AFLSDF_INV_57\);
    
    AFLSDF_INV_105 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_105\);
    
    \STAMP_0/spi/count[4]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[4]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_3\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[3]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_2_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[3]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_3_Z\, 
        CC => NET_CC_CONFIG113, P => NET_CC_CONFIG111, UB => 
        NET_CC_CONFIG112);
    
    AFLSDF_INV_63 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_63\);
    
    ResetAND_RNIMHJB : GB_NG
      port map(An => \AFLSDF_INV_49\, ENn => ADLIB_GND0, YNn => 
        OPEN, YSn => \ResetAND_RNIMHJB/U0_YNn_GSouth\);
    
    \MemorySynchronizer_0/resettimercounter_RNIV1O01[3]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_1978_i_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[3]\, C => 
        \MemorySynchronizer_0/un1_nreset_31_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[3]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_114\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[30]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[30]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[2]\, Y => 
        \MemorySynchronizer_0/N_1061\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[25]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[25]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[25]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[25]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[27]\ : SLE
      port map(D => \STAMP_0_data_frame[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[27]\);
    
    \MemorySynchronizer_0/dataReadyReset\ : SLE
      port map(D => \MemorySynchronizer_0/N_2068_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        ENABLE_MEMORY_LED_c, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => MemorySynchronizer_0_dataReadyReset);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4[10]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[10]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[10]\, C => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[10]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[14]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[14]\, B => 
        \sb_sb_0_STAMP_PWDATA[14]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[14]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_16\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[16]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[16]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_15\, S => 
        \MemorySynchronizer_0/temp_1[16]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_16\, CC => 
        NET_CC_CONFIG247, P => NET_CC_CONFIG245, UB => 
        NET_CC_CONFIG246);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_168\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data_2[8]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_591\, B => \STAMP_0/N_625\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_658\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_24\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[24]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_23_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[24]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_24_Z\, 
        CC => NET_CC_CONFIG176, P => NET_CC_CONFIG174, UB => 
        NET_CC_CONFIG175);
    
    \STAMP_0/un5_async_prescaler_count_cry_9\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[9]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_8_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_9_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_9_Z\, CC
         => NET_CC_CONFIG507, P => NET_CC_CONFIG505, UB => 
        NET_CC_CONFIG506);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_2\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[2]\, 
        B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_1_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_2_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_2_Z\, 
        CC => NET_CC_CONFIG633, P => NET_CC_CONFIG631, UB => 
        NET_CC_CONFIG632);
    
    AFLSDF_INV_30 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_30\);
    
    \STAMP_0/spi/count_cry[23]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[23]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[22]\, S => 
        \STAMP_0/spi/count_s[23]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[23]\, CC => NET_CC_CONFIG994, P
         => NET_CC_CONFIG992, UB => NET_CC_CONFIG993);
    
    \RXSM_LO_ibuf/U0/U_IOIN\ : IOIN_IB
      port map(YIN => \RXSM_LO_ibuf/U0/YIN\, E => ADLIB_GND0, Y
         => RXSM_LO_c);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_27_RNIUTGQ8\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[29]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[28]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[29]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[28]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[13]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[14]\, CC
         => NET_CC_CONFIG1159, P => NET_CC_CONFIG1157, UB => 
        NET_CC_CONFIG1158);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[31]\ : SLE
      port map(D => \STAMP_0_data_frame[31]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[31]\);
    
    \STAMP_0/un1_spi_rx_data_0[18]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[18]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[18]\, Y
         => \STAMP_0/N_601\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_2_0[20]\ : 
        CFG3
      generic map(INIT => x"0E")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\, 
        C => \MemorySynchronizer_0/SynchStatusReg_Z[23]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_2_0_Z[20]\);
    
    \STAMP_0/measurement_dms2[13]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[45]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[3]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_3_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_56\);
    
    AFLSDF_INV_92 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_40_Z\, Y => 
        \AFLSDF_INV_92\);
    
    \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa_1_i\ : 
        CFG4
      generic map(INIT => x"EAAA")

      port map(A => \MemorySynchronizer_0/N_2028_i\, B => 
        \MemorySynchronizer_0/N_2588\, C => 
        \MemorySynchronizer_0/APBState_Z[1]\, D => 
        \sb_sb_0_STAMP_PWDATA[30]\, Y => 
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa_1_i_Z\);
    
    \sb_sb_0/CoreAPB3_0/iPSELS_raw[0]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \sb_sb_0/STAMP_PADDRS[14]\, B => 
        \sb_sb_0/STAMP_PADDRS[13]\, C => 
        \sb_sb_0/CoreAPB3_0/iPSELS_raw_1_0_Z[0]\, D => 
        \sb_sb_0/STAMP_PADDRS[12]\, Y => sb_sb_0_STAMP_PSELx);
    
    AFLSDF_INV_66 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_46\, Y => 
        \AFLSDF_INV_66\);
    
    \MemorySynchronizer_0/TimeStampReg[25]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[25]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[25]\);
    
    \MemorySynchronizer_0/APBState_RNI199M[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \MemorySynchronizer_0/APBState_Z[0]\, B => 
        \MemorySynchronizer_0/APBState_Z[1]\, Y => 
        \MemorySynchronizer_0/N_301\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[26]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_26_S\, 
        Y => \MemorySynchronizer_0/N_1493\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_38\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[22]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_38_Z\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[20]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[20]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1071\, Y => 
        \MemorySynchronizer_0/N_1102\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_0_CC_0\ : 
        CC_CONFIG
      port map(CI => ADLIB_GND0, CO => CI_TO_CO293, P(0) => 
        NET_CC_CONFIG295, P(1) => NET_CC_CONFIG298, P(2) => 
        NET_CC_CONFIG301, P(3) => NET_CC_CONFIG304, P(4) => 
        NET_CC_CONFIG307, P(5) => NET_CC_CONFIG310, P(6) => 
        NET_CC_CONFIG313, P(7) => NET_CC_CONFIG316, P(8) => 
        NET_CC_CONFIG319, P(9) => NET_CC_CONFIG322, P(10) => 
        NET_CC_CONFIG325, P(11) => NET_CC_CONFIG328, UB(0) => 
        NET_CC_CONFIG296, UB(1) => NET_CC_CONFIG299, UB(2) => 
        NET_CC_CONFIG302, UB(3) => NET_CC_CONFIG305, UB(4) => 
        NET_CC_CONFIG308, UB(5) => NET_CC_CONFIG311, UB(6) => 
        NET_CC_CONFIG314, UB(7) => NET_CC_CONFIG317, UB(8) => 
        NET_CC_CONFIG320, UB(9) => NET_CC_CONFIG323, UB(10) => 
        NET_CC_CONFIG326, UB(11) => NET_CC_CONFIG329, CC(0) => 
        NET_CC_CONFIG297, CC(1) => NET_CC_CONFIG300, CC(2) => 
        NET_CC_CONFIG303, CC(3) => NET_CC_CONFIG306, CC(4) => 
        NET_CC_CONFIG309, CC(5) => NET_CC_CONFIG312, CC(6) => 
        NET_CC_CONFIG315, CC(7) => NET_CC_CONFIG318, CC(8) => 
        NET_CC_CONFIG321, CC(9) => NET_CC_CONFIG324, CC(10) => 
        NET_CC_CONFIG327, CC(11) => NET_CC_CONFIG330);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\);
    
    \MemorySynchronizer_0/ConfigReg[0]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[0]\);
    
    \STAMP_0/un1_pwdata[12]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[12]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => 
        \STAMP_0/un1_pwdata_Z[12]\);
    
    \STAMP_0/drdy_flank_detected_dms1_1_sqmuxa_1_i\ : CFG3
      generic map(INIT => x"FD")

      port map(A => stamp0_ready_dms1_c, B => 
        \STAMP_0/request_resync_0_sqmuxa\, C => 
        \STAMP_0/drdy_flank_detected_dms1_0_sqmuxa_1\, Y => 
        \STAMP_0/drdy_flank_detected_dms1_1_sqmuxa_1_i_Z\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_10\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_11\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_9_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[11]\, Y => OPEN, 
        FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_10_Z\, CC
         => NET_CC_CONFIG1053, P => NET_CC_CONFIG1051, UB => 
        NET_CC_CONFIG1052);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_27[10]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_2564\, C => 
        \MemorySynchronizer_0/N_271\, Y => 
        \MemorySynchronizer_0/N_2585\);
    
    \STAMP_0/measurement_temp[1]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[17]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[2]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[2]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1[30]\, Y => 
        \MemorySynchronizer_0/N_1089\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_13\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[13]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[13]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_12_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_13_Z\, CC => 
        NET_CC_CONFIG862, P => NET_CC_CONFIG860, UB => 
        NET_CC_CONFIG861);
    
    \MemorySynchronizer_0/un1_nreset_44_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_54_i_i_a2_Z\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_44_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_44_rs_Z\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[16]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[16]\, B => 
        \sb_sb_0_Memory_PRDATA[16]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[16]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[9]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[9]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[22]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[22]\);
    
    \STAMP_0/un1_spi_rx_data_0[29]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame[29]\, B => 
        \STAMP_0/config_Z[29]\, C => \sb_sb_0_STAMP_PADDR[8]\, Y
         => \STAMP_0/N_612\);
    
    AFLSDF_INV_44 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_42\, Y => 
        \AFLSDF_INV_44\);
    
    \STAMP_0/spi_tx_data_RNO[8]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[8]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_290_i\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_16\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_17\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_15_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[17]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_16_Z\, CC
         => NET_CC_CONFIG1071, P => NET_CC_CONFIG1069, UB => 
        NET_CC_CONFIG1070);
    
    \STAMP_0/spi/count_lm_0[17]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[17]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[17]\);
    
    
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa_i_1_i_a2_1\ : 
        CFG3
      generic map(INIT => x"02")

      port map(A => \MemorySynchronizer_0/APBState_Z[1]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, C => \sb_sb_0_STAMP_PADDR[5]\, 
        Y => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa_i_1_i_a2_1_Z\);
    
    \AND2_0_RNIKOS1/U0_RGB1\ : RGB_NG
      port map(An => \AND2_0_RNIKOS1/U0_YNn\, ENn => ADLIB_GND0, 
        YL => OPEN, YR => \AND2_0_RNIKOS1/U0_RGB1_YR\);
    
    \STAMP_0/un1_spi_rx_data[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0/N_651\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_5\, C => 
        \STAMP_0/spi_rx_data[1]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[1]\);
    
    \STAMP_0/component_state_RNO[5]\ : CFG4
      generic map(INIT => x"1113")

      port map(A => \STAMP_0/component_state_ns_0_i_a3_1_1_Z[0]\, 
        B => \STAMP_0/component_state_ns_0_i_0_0_Z[0]\, C => 
        \STAMP_0/N_109_i\, D => sb_sb_0_STAMP_PSELx, Y => 
        \STAMP_0/N_100_i\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[30]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[4]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[30]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[30]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[31]\ : CFG4
      generic map(INIT => x"1011")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[31]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[31]\, C => 
        \MemorySynchronizer_0/WaitingTimerValueReg_Z[31]\, D => 
        \MemorySynchronizer_0/N_1204_1\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[31]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_2_0[4]\ : 
        CFG4
      generic map(INIT => x"0020")

      port map(A => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, B
         => \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, C
         => \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[15]\, Y
         => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_2_0_Z[4]\);
    
    \STAMP_0/component_state_ns_0_0[2]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => \STAMP_0/spi_request_for_Z[0]\, B => 
        \STAMP_0/spi_request_for_Z[1]\, C => 
        \STAMP_0/component_state_ns_0_0_0_Z[2]\, D => 
        \STAMP_0/apb_spi_finished_0_sqmuxa_1\, Y => 
        \STAMP_0/component_state_ns[2]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[27]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[27]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[27]\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[27]\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[27]\);
    
    \STAMP_0/spi/count_lm_0[0]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => \STAMP_0/spi/count_Z[0]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[0]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[23]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[23]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[23]\, D
         => \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[23]\);
    
    \STAMP_0/async_prescaler_count[3]\ : SLE
      port map(D => \STAMP_0/un5_async_prescaler_count_cry_3_S\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[3]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[26]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_26_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[6]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/N_2588\, B => 
        \MemorySynchronizer_0/N_2597\, C => 
        \MemorySynchronizer_0/TimeStampReg_Z[4]\, D => 
        \MemorySynchronizer_0/ConfigReg_Z[4]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[4]\);
    
    \MemorySynchronizer_0/waitingtimercounter[27]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[27]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_38_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[27]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_34_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[2]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_34\);
    
    \MemorySynchronizer_0/un1_nreset_36_rs_RNI7NBL\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_43_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[29]\, C
         => \MemorySynchronizer_0/un1_nreset_36_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[29]\);
    
    \stamp0_ready_dms1_ibuf/U0/U_IOPAD\ : sdf_IOPAD_IN
      port map(PAD => stamp0_ready_dms1, Y => 
        \stamp0_ready_dms1_ibuf/U0/YIN1\);
    
    \MemorySynchronizer_0/TimeStampReg[15]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[15]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[15]\);
    
    \MemorySynchronizer_0/resynctimercounter[12]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1110\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[12]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_39\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_59_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_59\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_59_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_59_rs_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[28]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[28]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[28]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[4]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[28]\);
    
    \MemorySynchronizer_0/ConfigReg[17]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[17]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_3\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[3]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_2_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_3_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_3_Z\, CC
         => NET_CC_CONFIG734, P => NET_CC_CONFIG732, UB => 
        NET_CC_CONFIG733);
    
    AFLSDF_INV_75 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_75\);
    
    \STAMP_0/spi_tx_data[15]\ : SLE
      port map(D => \STAMP_0/N_268_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[15]\);
    
    \STAMP_0/un1_component_state_13_i_o2_RNO\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \STAMP_0/component_state_Z[5]\, B => 
        \STAMP_0/drdy_flank_detected_temp_Z\, C => 
        \STAMP_0/N_363\, D => \STAMP_0/N_158\, Y => 
        \STAMP_0/N_111_i\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[8]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[8]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[16]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[16]\, B => 
        \sb_sb_0_STAMP_PWDATA[16]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[16]\);
    
    \STAMP_0/component_state[1]\ : SLE
      port map(D => \STAMP_0/N_536_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/component_state_Z[1]\);
    
    \STAMP_0/un45_async_state_cry_3\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \STAMP_0/config_Z[27]\, B => 
        \STAMP_0_data_frame[6]\, C => ADLIB_GND0, D => ADLIB_GND0, 
        FCI => \STAMP_0/un45_async_state_cry_2_Z\, S => OPEN, Y
         => OPEN, FCO => \STAMP_0/un45_async_state_cry_3_Z\, CC
         => NET_CC_CONFIG525, P => NET_CC_CONFIG523, UB => 
        NET_CC_CONFIG524);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[24]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[24]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[23]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[24]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[24]\, CC
         => NET_CC_CONFIG78, P => NET_CC_CONFIG76, UB => 
        NET_CC_CONFIG77);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_60_set_RNIEJ5T\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_60_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[6]\, C
         => \MemorySynchronizer_0/un1_nreset_60_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[6]\);
    
    \MemorySynchronizer_0/TimeStampReg[3]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[3]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[3]\);
    
    \STAMP_0/un1_component_state_9_i_a3_1\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \STAMP_0/component_state_Z[4]\, B => 
        \STAMP_0/component_state_Z[2]\, C => 
        \STAMP_0/component_state_Z[0]\, D => \STAMP_0/N_160\, Y
         => \STAMP_0/un1_component_state_9_i_a3_1_Z\);
    
    AFLSDF_INV_18 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_54\, Y => 
        \AFLSDF_INV_18\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[21]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[21]\, B => 
        \sb_sb_0_Memory_PRDATA[21]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[21]\);
    
    \STAMP_0/un1_spi_rx_data_i_m2_1[30]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[62]\, B => 
        \STAMP_0/dummy_Z[30]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_220\);
    
    \nCS1_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => nCS1_c, E => ADLIB_VCC1, DOUT => 
        \nCS1_obuf/U0/DOUT1\, EOUT => \nCS1_obuf/U0/EOUT1\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a1_0\ : 
        CFG3
      generic map(INIT => x"02")

      port map(A => \MemorySynchronizer_0/APBState_Z[0]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, C => \sb_sb_0_STAMP_PADDR[6]\, 
        Y => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a1_0_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_268\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_YR\, C => ADLIB_VCC1, IPA
         => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CLK_BASE_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_27\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_28\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_26_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[28]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_27_Z\, CC
         => NET_CC_CONFIG1104, P => NET_CC_CONFIG1102, UB => 
        NET_CC_CONFIG1103);
    
    \STAMP_0/spi/count_lm_0[6]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[6]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[6]\);
    
    \STAMP_0/measurement_dms1[10]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[58]\);
    
    \STAMP_0/status_async_cycles_1_sqmuxa_1_i\ : CFG4
      generic map(INIT => x"5073")

      port map(A => \STAMP_0/un1_component_state_8_0_Z\, B => 
        \STAMP_0/async_state_Z[1]\, C => \STAMP_0/N_197\, D => 
        \STAMP_0/un1_async_prescaler_count\, Y => 
        \STAMP_0/status_async_cycles_1_sqmuxa_1_i_Z\);
    
    \MemorySynchronizer_0/PRDATA[8]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[8]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_5\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[5]\, 
        B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_4_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_5_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_5_Z\, 
        CC => NET_CC_CONFIG642, P => NET_CC_CONFIG640, UB => 
        NET_CC_CONFIG641);
    
    \STAMP_0/config[3]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[3]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[15]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[15]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[15]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[3]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[3]\, 
        B => \sb_sb_0_STAMP_PWDATA[3]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[3]\);
    
    \MemorySynchronizer_0/ConfigReg[1]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[1]\);
    
    \adc_clk_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => \sb_sb_0/CCC_0/GL1_INST/U0_RGB1_YR\, E => 
        ADLIB_VCC1, DOUT => \adc_clk_obuf/U0/DOUT1\, EOUT => 
        \adc_clk_obuf/U0/EOUT1\);
    
    \STAMP_0/apb_spi_finished_0_sqmuxa_1_0_a2\ : CFG3
      generic map(INIT => x"40")

      port map(A => \STAMP_0/spi_busy\, B => 
        \STAMP_0/component_state_Z[0]\, C => \STAMP_0/N_238\, Y
         => \STAMP_0/apb_spi_finished_0_sqmuxa_1\);
    
    \STAMP_0/spi/mosi_1\ : SLE
      port map(D => \STAMP_0/spi/tx_buffer_Z[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/mosi_1_1\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => mosi_1);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0[16]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[16]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[16]\, C => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[16]\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21[16]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10[28]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \MemorySynchronizer_0/N_2586\, B => 
        \MemorySynchronizer_0/N_2567\, Y => 
        \MemorySynchronizer_0/N_2588\);
    
    \MemorySynchronizer_0/MemorySyncState_RNI8R6JA[3]\ : CFG4
      generic map(INIT => x"8808")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => ENABLE_MEMORY_LED_c, C => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, D
         => \MemorySynchronizer_0/N_140_i_1\, Y => 
        \MemorySynchronizer_0/N_140_i\);
    
    \STAMP_0/un1_spi_rx_data_0[27]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame[27]\, B => 
        \STAMP_0/config_Z[27]\, C => \sb_sb_0_STAMP_PADDR[8]\, Y
         => \STAMP_0/N_610\);
    
    \STAMP_0/un1_new_avail_1_sqmuxa_3_i_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/N_238\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_333\);
    
    \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_1_0_a2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \STAMP_0/spi_request_for_Z[1]\, B => 
        \STAMP_0/spi_request_for_Z[0]\, C => 
        \STAMP_0/component_state_Z[0]\, D => \STAMP_0/N_331\, Y
         => \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14[28]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_18_0_Z[19]\, B
         => \MemorySynchronizer_0/N_271\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_Z[28]\, Y
         => \MemorySynchronizer_0/N_2596\);
    
    \STAMP_0/spi/un7_count_NE_13\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/spi/count_Z[24]\, B => 
        \STAMP_0/spi/count_Z[25]\, Y => 
        \STAMP_0/spi/un7_count_NE_13_Z\);
    
    \MemorySynchronizer_0/un1_nreset_27_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_55_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_27_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_27_rs_Z\);
    
    \MemorySynchronizer_0/TimeStampReg[8]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[8]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[8]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[29]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[29]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB0_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[29]\);
    
    \resetn_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => NN_1, E => ADLIB_VCC1, DOUT => 
        \resetn_obuf/U0/DOUT1\, EOUT => \resetn_obuf/U0/EOUT1\);
    
    \STAMP_0/un1_spi_rx_data[8]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_658\, C => \STAMP_0/spi_rx_data[8]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[8]\);
    
    \STAMP_0/spi/tx_buffer_RNO[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[15]\, B => 
        \STAMP_0/spi/tx_buffer_Z[14]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_120\);
    
    \STAMP_0/component_state_RNO[0]\ : CFG4
      generic map(INIT => x"0F08")

      port map(A => \STAMP_0/spi_busy\, B => 
        \STAMP_0/component_state_Z[1]\, C => \STAMP_0/N_331\, D
         => \STAMP_0/component_state_Z[0]\, Y => 
        \STAMP_0/N_487_i\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_17\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[17]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_16_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_17_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_17_Z\, 
        CC => NET_CC_CONFIG678, P => NET_CC_CONFIG676, UB => 
        NET_CC_CONFIG677);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_80\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_21_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_59_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_21_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_21_rs_Z\);
    
    \STAMP_0/delay_counter_cry[18]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[18]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[17]\, S
         => \STAMP_0/delay_counter_s[18]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[18]\, CC => NET_CC_CONFIG449, 
        P => NET_CC_CONFIG447, UB => NET_CC_CONFIG448);
    
    \STAMP_0/un68_paddr_1_0\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \sb_sb_0_STAMP_PADDR[8]\, B => 
        \STAMP_0/un52_paddr_5_Z\, C => \sb_sb_0_STAMP_PADDR[7]\, 
        D => \sb_sb_0_STAMP_PADDR[4]\, Y => 
        \STAMP_0/un68_paddr_1_0_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[9]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => \MemorySynchronizer_0/N_1182\, B => 
        \MemorySynchronizer_0/N_2575\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[9]\, D => 
        \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[9]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_46_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[26]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_46\);
    
    \STAMP_0/spi/count_cry[21]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[21]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[20]\, S => 
        \STAMP_0/spi/count_s[21]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[21]\, CC => NET_CC_CONFIG988, P
         => NET_CC_CONFIG986, UB => NET_CC_CONFIG987);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_2\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[2]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_1_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_2_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_2_Z\, CC
         => NET_CC_CONFIG731, P => NET_CC_CONFIG729, UB => 
        NET_CC_CONFIG730);
    
    \MemorySynchronizer_0/numberofnewavails_RNI0D491[0]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[0]\, 
        B => \MemorySynchronizer_0/N_140_2\, C => 
        \MemorySynchronizer_0/numberofnewavails_Z[2]\, D => 
        \MemorySynchronizer_0/numberofnewavails_Z[1]\, Y => 
        \MemorySynchronizer_0/N_2321\);
    
    AFLSDF_INV_3 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_41_Z\, Y => 
        \AFLSDF_INV_3\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_170\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_38_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_50\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_38_set_Z\);
    
    \STAMP_0/un45_async_state_cry_0\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \STAMP_0/config_Z[24]\, B => 
        \STAMP_0_data_frame[3]\, C => ADLIB_GND0, D => ADLIB_GND0, 
        FCI => ADLIB_GND0, S => OPEN, Y => OPEN, FCO => 
        \STAMP_0/un45_async_state_cry_0_Z\, CC => 
        NET_CC_CONFIG516, P => NET_CC_CONFIG514, UB => 
        NET_CC_CONFIG515);
    
    \ENABLE_MEMORY_LED_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \ENABLE_MEMORY_LED_obuf/U0/EOUT1\, Y => 
        \ENABLE_MEMORY_LED_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[22]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_22\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[22]\, 
        C => \MemorySynchronizer_0/N_1501\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[22]\);
    
    \MemorySynchronizer_0/un1_nreset_47_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[16]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_47_i\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[0]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_0\);
    
    \RXSM_LO_ibuf/U0/U_IOPAD\ : sdf_IOPAD_IN
      port map(PAD => RXSM_LO, Y => \RXSM_LO_ibuf/U0/YIN1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[18]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[18]\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2564\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1437\);
    
    \MemorySynchronizer_0/un1_nreset_26_rs_RNI1C3J\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_51_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[25]\, C
         => \MemorySynchronizer_0/un1_nreset_26_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[25]\);
    
    \STAMP_0/un1_component_state_13_i_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \STAMP_0/component_state_Z[4]\, B => 
        \STAMP_0/component_state_Z[1]\, C => \STAMP_0/N_155\, D
         => \STAMP_0/N_156\, Y => \STAMP_0/N_337\);
    
    \MemorySynchronizer_0/SynchStatusReg2[25]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[25]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[25]\);
    
    \MemorySynchronizer_0/resynctimercounter[18]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1104\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[18]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[5]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[5]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[4]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[5]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[5]\, CC
         => NET_CC_CONFIG21, P => NET_CC_CONFIG19, UB => 
        NET_CC_CONFIG20);
    
    \MemorySynchronizer_0/un1_nreset_3_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/N_21_i\, EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_3_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_3_rs_Z\);
    
    \STAMP_0/spi/rx_data[0]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB0_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[0]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[10]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_10\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[10]\, 
        C => \MemorySynchronizer_0/N_2434\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[10]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_52_set_RNIVCEF\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_52_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[14]\, C
         => \MemorySynchronizer_0/un1_nreset_52_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[14]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_58\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[4]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_ResetTimerValueReg_58_Z\);
    
    \STAMP_0/spi_tx_data[5]\ : SLE
      port map(D => \STAMP_0/N_293_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[5]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[21]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[21]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[11]\, Y
         => \MemorySynchronizer_0/N_1070\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_233\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[29]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[29]\, B => 
        \sb_sb_0_STAMP_PWDATA[29]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[29]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[15]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[15]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1076\, Y => 
        \MemorySynchronizer_0/N_1107\);
    
    \MemorySynchronizer_0/resettimercounter_RNIF1AQ[4]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_58_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[4]\, C => 
        \MemorySynchronizer_0/un1_nreset_30_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[4]\);
    
    \STAMP_0/spi_tx_data[13]\ : SLE
      port map(D => \STAMP_0/N_266_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[13]\);
    
    \STAMP_0/spi/count[30]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[30]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB12_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[30]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[9]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[9]\, 
        B => \sb_sb_0_STAMP_PWDATA[9]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[9]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_3\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[3]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[3]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_2\, S => 
        \MemorySynchronizer_0/temp_1[3]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_3\, CC => 
        NET_CC_CONFIG208, P => NET_CC_CONFIG206, UB => 
        NET_CC_CONFIG207);
    
    \MemorySynchronizer_0/un1_nreset_9\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[24]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_9_i\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_19\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[19]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_18_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_19_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_19_Z\, 
        CC => NET_CC_CONFIG684, P => NET_CC_CONFIG682, UB => 
        NET_CC_CONFIG683);
    
    \STAMP_0/spi_tx_data_RNO[9]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[9]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_289_i\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[11]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[11]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[11]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[22]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[22]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[22]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[22]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[6]\ : SLE
      port map(D => \STAMP_0_data_frame[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[6]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[10]\ : SLE
      port map(D => \STAMP_0_data_frame[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[10]\);
    
    \STAMP_0/measurement_dms2[15]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[47]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[4]\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[4]\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[4]\, C => 
        \MemorySynchronizer_0/N_2593\, D => 
        \MemorySynchronizer_0/N_1260\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[4]\);
    
    \STAMP_0/spi/count[9]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[9]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[7]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[7]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[31]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[31]\, B => 
        \sb_sb_0_Memory_PRDATA[31]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[31]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_0_CC_2\ : CC_CONFIG
      port map(CI => CI_TO_CO820, CO => OPEN, P(0) => 
        NET_CC_CONFIG893, P(1) => NET_CC_CONFIG896, P(2) => 
        NET_CC_CONFIG899, P(3) => NET_CC_CONFIG902, P(4) => 
        NET_CC_CONFIG905, P(5) => NET_CC_CONFIG908, P(6) => 
        NET_CC_CONFIG911, P(7) => NET_CC_CONFIG914, P(8) => 
        NET_CC_CONFIG917, P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, 
        P(11) => ADLIB_VCC1, UB(0) => NET_CC_CONFIG894, UB(1) => 
        NET_CC_CONFIG897, UB(2) => NET_CC_CONFIG900, UB(3) => 
        NET_CC_CONFIG903, UB(4) => NET_CC_CONFIG906, UB(5) => 
        NET_CC_CONFIG909, UB(6) => NET_CC_CONFIG912, UB(7) => 
        NET_CC_CONFIG915, UB(8) => NET_CC_CONFIG918, UB(9) => 
        ADLIB_VCC1, UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, 
        CC(0) => NET_CC_CONFIG895, CC(1) => NET_CC_CONFIG898, 
        CC(2) => NET_CC_CONFIG901, CC(3) => NET_CC_CONFIG904, 
        CC(4) => NET_CC_CONFIG907, CC(5) => NET_CC_CONFIG910, 
        CC(6) => NET_CC_CONFIG913, CC(7) => NET_CC_CONFIG916, 
        CC(8) => NET_CC_CONFIG919, CC(9) => nc395, CC(10) => 
        nc280, CC(11) => nc125);
    
    \STAMP_0/un1_new_avail_1_sqmuxa_3_i_0\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/un1_new_avail_0_sqmuxa_1\, B => 
        \STAMP_0/N_333\, Y => 
        \STAMP_0/un1_new_avail_1_sqmuxa_3_i_0_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[3]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_56\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[3]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[3]\, D
         => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[3]\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_0\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/CLK0_net\, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/PSEL_net\, IPC => OPEN);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_16\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[22]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[21]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[19]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[15]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_16_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[25]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[25]\, B => 
        \sb_sb_0_STAMP_PWDATA[25]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[25]\);
    
    \STAMP_0/status_async_cycles_s_388_CC_0\ : CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => OPEN, P(0) => ADLIB_VCC1, 
        P(1) => ADLIB_VCC1, P(2) => ADLIB_GND0, P(3) => 
        NET_CC_CONFIG587, P(4) => NET_CC_CONFIG590, P(5) => 
        NET_CC_CONFIG593, P(6) => NET_CC_CONFIG596, P(7) => 
        NET_CC_CONFIG599, P(8) => NET_CC_CONFIG602, P(9) => 
        ADLIB_VCC1, P(10) => ADLIB_VCC1, P(11) => ADLIB_VCC1, 
        UB(0) => ADLIB_VCC1, UB(1) => ADLIB_VCC1, UB(2) => 
        ADLIB_GND0, UB(3) => NET_CC_CONFIG588, UB(4) => 
        NET_CC_CONFIG591, UB(5) => NET_CC_CONFIG594, UB(6) => 
        NET_CC_CONFIG597, UB(7) => NET_CC_CONFIG600, UB(8) => 
        NET_CC_CONFIG603, UB(9) => ADLIB_VCC1, UB(10) => 
        ADLIB_VCC1, UB(11) => ADLIB_VCC1, CC(0) => nc211, CC(1)
         => nc73, CC(2) => nc107, CC(3) => NET_CC_CONFIG589, 
        CC(4) => NET_CC_CONFIG592, CC(5) => NET_CC_CONFIG595, 
        CC(6) => NET_CC_CONFIG598, CC(7) => NET_CC_CONFIG601, 
        CC(8) => NET_CC_CONFIG604, CC(9) => nc408, CC(10) => 
        nc329, CC(11) => nc66);
    
    \MemorySynchronizer_0/ConfigReg_0_0_a3_0_a2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \MemorySynchronizer_0/APBState_Z[0]\, B => 
        \MemorySynchronizer_0/APBState_Z[1]\, C => 
        \MemorySynchronizer_0/N_2586\, D => 
        \MemorySynchronizer_0/N_2567\, Y => 
        \MemorySynchronizer_0/ConfigReg_0\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_13_RNIBIFT7\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[15]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[14]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[15]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[14]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[6]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[7]\, CC
         => NET_CC_CONFIG1138, P => NET_CC_CONFIG1136, UB => 
        NET_CC_CONFIG1137);
    
    \STAMP_0/async_state_0_sqmuxa_1_1\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \STAMP_0/apb_is_reset_Z\, B => 
        \STAMP_0/async_state_Z[0]\, C => 
        \STAMP_0/async_state_Z[1]\, D => 
        \STAMP_0/component_state_Z[2]\, Y => 
        \STAMP_0/async_state_0_sqmuxa_1_1_Z\);
    
    \STAMP_0/spi/count_cry[5]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[5]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[4]\, S => 
        \STAMP_0/spi/count_s[5]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[5]\, CC => NET_CC_CONFIG940, P
         => NET_CC_CONFIG938, UB => NET_CC_CONFIG939);
    
    \stamp0_spi_miso_ibuf/U0/U_IOPAD\ : sdf_IOPAD_IN
      port map(PAD => stamp0_spi_miso, Y => 
        \stamp0_spi_miso_ibuf/U0/YIN1\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[7]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[7]\, B => 
        \sb_sb_0_Memory_PRDATA[7]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7]\);
    
    \STAMP_0/measurement_dms1[2]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[50]\);
    
    \STAMP_0/drdy_flank_detected_dms2\ : SLE
      port map(D => \STAMP_0/stamp0_ready_dms2_c_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/drdy_flank_detected_dms2_1_sqmuxa_2_i_Z\, ALn
         => \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/drdy_flank_detected_dms2_Z\);
    
    \MemorySynchronizer_0/PRDATA[31]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[31]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[31]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_132\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[17]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[17]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[10]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[10]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[10]\);
    
    \STAMP_0/un1_component_state_14_i_0\ : CFG4
      generic map(INIT => x"AE00")

      port map(A => \STAMP_0/N_364\, B => \STAMP_0/N_248_2\, C
         => \STAMP_0/spi_request_for_Z[0]\, D => \STAMP_0/N_165\, 
        Y => \STAMP_0/un1_component_state_14_i_0_Z\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_31_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_51\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_31_set_Z\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_1\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[1]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_0_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[31]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_1_Z\, CC
         => NET_CC_CONFIG300, P => NET_CC_CONFIG298, UB => 
        NET_CC_CONFIG299);
    
    \MemorySynchronizer_0/PRDATA[5]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[5]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[5]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[17]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_17_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[15]\);
    
    \STAMP_0/request_resync_1_sqmuxa_1\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \STAMP_0/async_state_Z[1]\, B => 
        \STAMP_0/async_state_Z[0]\, C => 
        \STAMP_0/un1_async_prescaler_count\, D => 
        \STAMP_0/un45_async_state_cry_5_Z\, Y => 
        \STAMP_0/request_resync_1_sqmuxa_1_Z\);
    
    \STAMP_0/spi/sclk_buffer_RNO\ : CFG4
      generic map(INIT => x"2788")

      port map(A => \STAMP_0/spi/state_Z[0]\, B => 
        \STAMP_0/spi/sclk_buffer_0_sqmuxa\, C => \STAMP_0/enable\, 
        D => stamp0_spi_clock_c, Y => \STAMP_0/spi/N_20_i\);
    
    \MemorySynchronizer_0/resynctimercounter[4]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1118\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[4]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_58_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_52\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_58_set_Z\);
    
    \STAMP_0/delay_counter_lm_0[10]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[10]\, Y => 
        \STAMP_0/delay_counter_lm[10]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[26]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[26]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[6]\, Y => 
        \MemorySynchronizer_0/N_1065\);
    
    \STAMP_0/delay_counter[2]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[2]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS_1[1]\ : CFG4
      generic map(INIT => x"40C0")

      port map(A => \sb_sb_0/STAMP_PADDRS[14]\, B => 
        \sb_sb_0/STAMP_PADDRS[13]\, C => 
        \sb_sb_0/CoreAPB3_0/iPSELS_raw_1_0_Z[0]\, D => 
        \sb_sb_0/STAMP_PADDRS[12]\, Y => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS[1]\);
    
    \STAMP_0/measurement_temp[8]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[24]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[7]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \MemorySynchronizer_0/N_2585\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[7]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[7]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[7]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[15]\ : SLE
      port map(D => \STAMP_0_data_frame[47]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[15]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[14]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[14]\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/N_2323\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[14]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[14]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_235\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_6[1]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[1]\, 
        B => \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2567\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1177\);
    
    \STAMP_0/spi_request_for_2_sqmuxa_0_o2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/drdy_flank_detected_dms1_Z\, B => 
        \STAMP_0/drdy_flank_detected_dms2_Z\, Y => 
        \STAMP_0/N_158\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_140\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_EV_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv[11]\ : CFG4
      generic map(INIT => x"EECE")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[13]\, 
        B => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_1_Z[11]\, C
         => \MemorySynchronizer_0/N_6\, D => 
        \MemorySynchronizer_0/N_1512\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168[11]\);
    
    \LED_HEARTBEAT_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \LED_HEARTBEAT_obuf/U0/EOUT1\, Y => 
        \LED_HEARTBEAT_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/ConfigReg[4]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[4]\);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_22\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[14]\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[12]\, C => 
        \MemorySynchronizer_0/waitingtimercounter_Z[11]\, D => 
        \MemorySynchronizer_0/waitingtimercounter_Z[8]\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_22_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[2]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[2]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[1]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[2]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[2]\, CC
         => NET_CC_CONFIG12, P => NET_CC_CONFIG10, UB => 
        NET_CC_CONFIG11);
    
    \stamp0_spi_dms1_cs_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \stamp0_spi_dms1_cs_obuf/U0/EOUT1\, Y => 
        \stamp0_spi_dms1_cs_obuf/U0/EOUT\);
    
    AFLSDF_INV_71 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_71\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_16\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[16]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_15_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[16]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_16_Z\, CC
         => NET_CC_CONFIG345, P => NET_CC_CONFIG343, UB => 
        NET_CC_CONFIG344);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[17]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[17]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[15]\, Y
         => \MemorySynchronizer_0/N_1074\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[27]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[27]\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/N_2323\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[27]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[27]\);
    
    \MemorySynchronizer_0/waitingtimercounter_RNI1P0Q[12]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_54_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[12]\, C
         => \MemorySynchronizer_0/un1_nreset_54_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[12]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_4_0[20]\ : 
        CFG3
      generic map(INIT => x"0E")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\, 
        C => \MemorySynchronizer_0/SynchStatusReg_Z[26]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_4_0_Z[20]\);
    
    \STAMP_0/spi/count_lm_0[21]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[21]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[21]\);
    
    \MemorySynchronizer_0/TimeStampGen/un1_prescaler_ac0_1\ : 
        CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/enableTimestampGen_Z\, 
        B => \MemorySynchronizer_0/TimeStampGen/prescaler_Z[1]\, 
        C => \MemorySynchronizer_0/TimeStampGen/prescaler_Z[0]\, 
        Y => \MemorySynchronizer_0/TimeStampGen/un1_prescaler_c2\);
    
    \STAMP_0/config[26]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[26]\);
    
    \stamp0_ready_temp_ibuf/U0/U_IOIN\ : IOIN_IB
      port map(YIN => \stamp0_ready_temp_ibuf/U0/YIN\, E => 
        ADLIB_GND0, Y => stamp0_ready_temp_c);
    
    \MemorySynchronizer_0/un1_nreset_15_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[18]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_15_i\);
    
    AFLSDF_INV_54 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_54\);
    
    \STAMP_0/delay_counter_lm_0[11]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[11]\, Y => 
        \STAMP_0/delay_counter_lm[11]\);
    
    \MemorySynchronizer_0/resettimercounter[22]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_11_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[22]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[27]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[1]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[27]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[27]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[23]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_23\);
    
    \MemorySynchronizer_0/N_1979_i_set_RNIOTBQ\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_1979_i_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[15]\, C => 
        \MemorySynchronizer_0/un1_nreset_18_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[15]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_18_0[19]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_18_0_Z[19]\);
    
    \MemorySynchronizer_0/resettimercounter[17]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_16_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[17]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0[8]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[8]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[8]\, C => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[8]\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21[8]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[28]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_28\);
    
    \STAMP_0/spi/count_lm_0[3]\ : CFG4
      generic map(INIT => x"D8CC")

      port map(A => \STAMP_0/spi/un7_count_NE_i\, B => 
        \STAMP_0/spi/count_0_sqmuxa\, C => 
        \STAMP_0/spi/count_s[3]\, D => \STAMP_0/spi/state_Z[0]\, 
        Y => \STAMP_0/spi/count_lm[3]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_42\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[18]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_42_Z\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_8\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[8]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_7_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[24]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_8_Z\, CC
         => NET_CC_CONFIG321, P => NET_CC_CONFIG319, UB => 
        NET_CC_CONFIG320);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_0_CC_2\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO1020, CO => OPEN, P(0) => 
        NET_CC_CONFIG1084, P(1) => NET_CC_CONFIG1087, P(2) => 
        NET_CC_CONFIG1090, P(3) => NET_CC_CONFIG1093, P(4) => 
        NET_CC_CONFIG1096, P(5) => NET_CC_CONFIG1099, P(6) => 
        NET_CC_CONFIG1102, P(7) => NET_CC_CONFIG1105, P(8) => 
        NET_CC_CONFIG1108, P(9) => NET_CC_CONFIG1111, P(10) => 
        ADLIB_VCC1, P(11) => ADLIB_VCC1, UB(0) => 
        NET_CC_CONFIG1085, UB(1) => NET_CC_CONFIG1088, UB(2) => 
        NET_CC_CONFIG1091, UB(3) => NET_CC_CONFIG1094, UB(4) => 
        NET_CC_CONFIG1097, UB(5) => NET_CC_CONFIG1100, UB(6) => 
        NET_CC_CONFIG1103, UB(7) => NET_CC_CONFIG1106, UB(8) => 
        NET_CC_CONFIG1109, UB(9) => NET_CC_CONFIG1112, UB(10) => 
        ADLIB_VCC1, UB(11) => ADLIB_VCC1, CC(0) => 
        NET_CC_CONFIG1086, CC(1) => NET_CC_CONFIG1089, CC(2) => 
        NET_CC_CONFIG1092, CC(3) => NET_CC_CONFIG1095, CC(4) => 
        NET_CC_CONFIG1098, CC(5) => NET_CC_CONFIG1101, CC(6) => 
        NET_CC_CONFIG1104, CC(7) => NET_CC_CONFIG1107, CC(8) => 
        NET_CC_CONFIG1110, CC(9) => NET_CC_CONFIG1113, CC(10) => 
        nc83, CC(11) => nc9);
    
    
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_3_i_0_a2_1_RNITIUG1\ : 
        CFG4
      generic map(INIT => x"7333")

      port map(A => \MemorySynchronizer_0/APBState_Z[0]\, B => 
        \MemorySynchronizer_0/N_301\, C => 
        \MemorySynchronizer_0/N_2567\, D => 
        \MemorySynchronizer_0/N_2586\, Y => 
        \MemorySynchronizer_0/un1_APBState_i\);
    
    \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_4\ : 
        CFG4
      generic map(INIT => x"E000")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[0]\, 
        B => \MemorySynchronizer_0/MemorySyncState_Z[2]\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_29_Z\, 
        D => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_30_Z\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_4_Z\);
    
    \STAMP_0/spi/tx_buffer_RNO[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[11]\, B => 
        \STAMP_0/spi/tx_buffer_Z[10]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_124\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_3\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[3]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_2_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[29]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_3_Z\, CC
         => NET_CC_CONFIG306, P => NET_CC_CONFIG304, UB => 
        NET_CC_CONFIG305);
    
    \STAMP_0/delay_counter_RNIMTFR[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \STAMP_0/delay_counter_Z[7]\, B => 
        \STAMP_0/delay_counter_Z[6]\, C => 
        \STAMP_0/delay_counter_Z[5]\, D => 
        \STAMP_0/delay_counter_Z[4]\, Y => 
        \STAMP_0/N_517_i_0_a2_19\);
    
    \MemorySynchronizer_0/TimeStampReg[27]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[27]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[27]\);
    
    \STAMP_0/un1_component_state_13_i_o2_0\ : CFG3
      generic map(INIT => x"57")

      port map(A => \STAMP_0/component_state_Z[2]\, B => 
        sb_sb_0_STAMP_PENABLE, C => \STAMP_0/apb_is_atomic_Z\, Y
         => \STAMP_0/N_156\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_187\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/ResetTimerValueReg[28]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[28]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[2]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_2\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[2]\, 
        C => \MemorySynchronizer_0/N_1565\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[2]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[4]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[4]\, C => 
        \MemorySynchronizer_0/N_2596\, D => 
        \MemorySynchronizer_0/N_2595\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[4]\);
    
    \nCS2_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => nCS2, D => \nCS2_obuf/U0/DOUT\, E => 
        \nCS2_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_17\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[17]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_16_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[15]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_17_Z\, CC
         => NET_CC_CONFIG348, P => NET_CC_CONFIG346, UB => 
        NET_CC_CONFIG347);
    
    AFLSDF_INV_48 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_33_Z\, Y => 
        \AFLSDF_INV_48\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[13]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[13]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_15\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_16\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_14_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[16]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_15_Z\, CC
         => NET_CC_CONFIG1068, P => NET_CC_CONFIG1066, UB => 
        NET_CC_CONFIG1067);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_4\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[4]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[4]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_3\, S => 
        \MemorySynchronizer_0/temp_1[4]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_4\, CC => 
        NET_CC_CONFIG211, P => NET_CC_CONFIG209, UB => 
        NET_CC_CONFIG210);
    
    \STAMP_0/spi/clk_toggles_cry[4]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/spi/clk_toggles_Z[4]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/spi/clk_toggles_cry_Z[3]\, S
         => \STAMP_0/spi/clk_toggles_s[4]\, Y => OPEN, FCO => 
        \STAMP_0/spi/clk_toggles_cry_Z[4]\, CC => 
        NET_CC_CONFIG619, P => NET_CC_CONFIG617, UB => 
        NET_CC_CONFIG618);
    
    \MemorySynchronizer_0/ResetTimerValueReg[24]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[24]\);
    
    \MemorySynchronizer_0/PRDATA[17]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[17]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[17]\);
    
    \MemorySynchronizer_0/waitingtimercounter_RNI4K901[16]\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_33_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[16]\, C
         => \MemorySynchronizer_0/un1_nreset_47_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[16]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_32\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_20_rs_RNI9F351\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_47_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[0]\, C
         => \MemorySynchronizer_0/un1_nreset_20_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[0]\);
    
    \STAMP_0/spi/clk_toggles_cry[3]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/spi/clk_toggles_Z[3]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/spi/clk_toggles_cry_Z[2]\, S
         => \STAMP_0/spi/clk_toggles_s[3]\, Y => OPEN, FCO => 
        \STAMP_0/spi/clk_toggles_cry_Z[3]\, CC => 
        NET_CC_CONFIG616, P => NET_CC_CONFIG614, UB => 
        NET_CC_CONFIG615);
    
    \STAMP_0/un1_spi_rx_data_0[9]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[9]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[9]\, Y
         => \STAMP_0/N_592\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_55_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[11]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_55\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[3]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_3\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_0_Z[3]\, 
        C => \MemorySynchronizer_0/N_1209\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[3]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_RNO_0[5]\ : 
        CFG4
      generic map(INIT => x"0C05")

      port map(A => STAMP_0_new_avail, B => 
        \MemorySynchronizer_0/SynchStatusReg_Z[7]\, C => 
        \MemorySynchronizer_0/N_6\, D => 
        \MemorySynchronizer_0/SynchStatusReg_N_7\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_82_m[5]\);
    
    \MemorySynchronizer_0/resynctimercounter[16]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1106\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[16]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_14\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[14]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_13_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[14]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_14_Z\, 
        CC => NET_CC_CONFIG146, P => NET_CC_CONFIG144, UB => 
        NET_CC_CONFIG145);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[25]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_25\);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB9\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_21\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[20]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[13]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[8]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[6]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_21_Z\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[5]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[5]\);
    
    \MemorySynchronizer_0/waitingtimercounter[15]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[15]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_51_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[15]\);
    
    \MemorySynchronizer_0/un1_nreset_45_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_34\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_45_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_45_rs_Z\);
    
    \STAMP_0/un1_spi_rx_data[7]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_657\, C => \STAMP_0/spi_rx_data[7]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[7]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_45_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_53\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_45_set_Z\);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_22\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[30]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[28]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[16]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[1]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_22_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[7]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_7_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_64\);
    
    \MemorySynchronizer_0/un1_nreset_62_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[20]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_62_i\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_23\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[23]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_22_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_23_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_23_Z\, CC
         => NET_CC_CONFIG794, P => NET_CC_CONFIG792, UB => 
        NET_CC_CONFIG793);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_34_RNO[20]\ : 
        CFG4
      generic map(INIT => x"2A0A")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => \MemorySynchronizer_0/g0_0_1\, C => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, D
         => \MemorySynchronizer_0/N_140_2\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_34_1[20]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[5]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[5]\);
    
    \MemorySynchronizer_0/TimeStampReg[17]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[17]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[17]\);
    
    \STAMP_0/un1_component_state_8_0\ : CFG3
      generic map(INIT => x"27")

      port map(A => \STAMP_0/component_state_Z[5]\, B => 
        \STAMP_0/config_Z[31]\, C => 
        \STAMP_0/component_state_Z[0]\, Y => 
        \STAMP_0/un1_component_state_8_0_Z\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[25]\ : SLE
      port map(D => \STAMP_0_data_frame[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[25]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_13\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[18]\, B
         => ADLIB_VCC1, C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18]\, 
        IPB => OPEN, IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_206\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_23_RNIQ97I8\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[25]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[24]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[25]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[24]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[11]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[12]\, CC
         => NET_CC_CONFIG1153, P => NET_CC_CONFIG1151, UB => 
        NET_CC_CONFIG1152);
    
    \STAMP_0/component_state_ns_0[3]\ : CFG4
      generic map(INIT => x"8F0F")

      port map(A => \STAMP_0/component_state_Z[3]\, B => 
        \STAMP_0/apb_spi_finished_Z\, C => 
        \STAMP_0/component_state_ns_0_1_Z[3]\, D => 
        \STAMP_0/un27_paddr_i_0\, Y => 
        \STAMP_0/component_state_ns[3]\);
    
    \STAMP_0/un1_spi_rx_data_2[12]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_595\, B => \STAMP_0/N_629\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_662\);
    
    \STAMP_0/dummy[15]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_54\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[15]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[1]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_1\);
    
    \MemorySynchronizer_0/un1_nreset_33_0_a3_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[1]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_33_i\);
    
    \MemorySynchronizer_0/MemorySyncState[5]\ : SLE
      port map(D => \MemorySynchronizer_0/MemorySyncState_ns[0]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, 
        EN => ENABLE_MEMORY_LED_c, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/MemorySyncState_Z[5]\);
    
    AFLSDF_INV_110 : INV_BA
      port map(A => \sb_sb_0/CCC_0/GL0_net\, Y => 
        \AFLSDF_INV_110\);
    
    \STAMP_0/un1_spi_rx_data_sn_m4_0_a3\ : CFG2
      generic map(INIT => x"1")

      port map(A => \sb_sb_0_STAMP_PADDR[8]\, B => 
        \sb_sb_0_STAMP_PADDR[9]\, Y => 
        \STAMP_0/un1_spi_rx_data_sn_N_5\);
    
    \MemorySynchronizer_0/SynchStatusReg2[2]\ : SLE
      port map(D => \MemorySynchronizer_0/temp_1[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[2]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[6]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[6]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1085\, Y => 
        \MemorySynchronizer_0/N_1116\);
    
    \nCS2_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \nCS2_obuf/U0/EOUT1\, Y => 
        \nCS2_obuf/U0/EOUT\);
    
    AFLSDF_INV_10 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_38_Z\, Y => 
        \AFLSDF_INV_10\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_87\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[29]\, B => 
        \MemorySynchronizer_0/un104_in_enable_28\, C => 
        \MemorySynchronizer_0/un104_in_enable_29\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[28]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[13]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[14]\, CC
         => NET_CC_CONFIG580, P => NET_CC_CONFIG578, UB => 
        NET_CC_CONFIG579);
    
    \STAMP_0/spi/count_cry[4]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[4]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[3]\, S => 
        \STAMP_0/spi/count_s[4]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[4]\, CC => NET_CC_CONFIG937, P
         => NET_CC_CONFIG935, UB => NET_CC_CONFIG936);
    
    \STAMP_0/status_async_cycles_cry[4]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0_data_frame[7]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/status_async_cycles_cry_Z[3]\, S => 
        \STAMP_0/status_async_cycles_s[4]\, Y => OPEN, FCO => 
        \STAMP_0/status_async_cycles_cry_Z[4]\, CC => 
        NET_CC_CONFIG601, P => NET_CC_CONFIG599, UB => 
        NET_CC_CONFIG600);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_81\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22]\, 
        IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data_2[2]\ : CFG4
      generic map(INIT => x"D155")

      port map(A => \STAMP_0/un1_spi_rx_data_2_1_0_Z[2]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/dummy_Z[2]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_652\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO[25]\ : CFG4
      generic map(INIT => x"050D")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_3_0_Z[20]\, 
        B => \MemorySynchronizer_0/N_2321\, C => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, D => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\, 
        Y => \MemorySynchronizer_0/N_2033_i\);
    
    \STAMP_0/spi/count_cry[19]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[19]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[18]\, S => 
        \STAMP_0/spi/count_s[19]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[19]\, CC => NET_CC_CONFIG982, P
         => NET_CC_CONFIG980, UB => NET_CC_CONFIG981);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[16]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[16]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[16]\, C => 
        \MemorySynchronizer_0/N_2596\, D => 
        \MemorySynchronizer_0/N_2595\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[16]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[15]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[15]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[15]\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[15]\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[15]\);
    
    \STAMP_0/delay_counter_cry[16]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[16]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[15]\, S
         => \STAMP_0/delay_counter_s[16]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[16]\, CC => NET_CC_CONFIG443, 
        P => NET_CC_CONFIG441, UB => NET_CC_CONFIG442);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_o2[31]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => \MemorySynchronizer_0/N_2561\, B => 
        \MemorySynchronizer_0/N_2567\, C => 
        \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/N_1123\);
    
    AFLSDF_INV_112 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_112\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_16[20]\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[26]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[25]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[24]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[23]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_16_Z[20]\);
    
    \STAMP_0/spi/assert_data_5_iv_0_a2_0\ : CFG3
      generic map(INIT => x"40")

      port map(A => \STAMP_0/spi/assert_data_Z\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => \STAMP_0/spi/N_63\);
    
    \STAMP_0/delay_counter[6]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[6]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[8]\ : SLE
      port map(D => \STAMP_0_data_frame[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[8]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_202\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[29]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[29]\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2564\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1403\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_22\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/N_1088\, B => 
        \MemorySynchronizer_0/N_1086\, C => 
        \MemorySynchronizer_0/N_1071\, D => 
        \MemorySynchronizer_0/N_1069\, Y => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_22_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[13]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_13\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[13]\, 
        C => \MemorySynchronizer_0/N_1525\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[13]\);
    
    \LED_HEARTBEAT_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \LED_HEARTBEAT_obuf/U0/DOUT1\, Y => 
        \LED_HEARTBEAT_obuf/U0/DOUT\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_35\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_1_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_49\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_1_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_1_rs_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[26]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[26]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[28]\, C => 
        \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_1182\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[26]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_131\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[28]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[28]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[28]\, C => 
        \MemorySynchronizer_0/N_2596\, D => 
        \MemorySynchronizer_0/N_2595\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[28]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[25]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[25]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[25]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[7]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[25]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_25\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un104_in_enable_25\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[25]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_24_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_25_Z\, CC => 
        NET_CC_CONFIG898, P => NET_CC_CONFIG896, UB => 
        NET_CC_CONFIG897);
    
    AFLSDF_INV_108 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_55_Z\, Y => 
        \AFLSDF_INV_108\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_23\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[23]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_22_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[9]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_23_Z\, CC
         => NET_CC_CONFIG366, P => NET_CC_CONFIG364, UB => 
        NET_CC_CONFIG365);
    
    \STAMP_0/PRDATA[15]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[15]\);
    
    \STAMP_0/delay_counter_cry[3]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[3]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/delay_counter_cry_Z[2]\, S => 
        \STAMP_0/delay_counter_s[3]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[3]\, CC => NET_CC_CONFIG404, 
        P => NET_CC_CONFIG402, UB => NET_CC_CONFIG403);
    
    \STAMP_0/spi/tx_buffer[4]\ : SLE
      port map(D => \STAMP_0/spi/N_134\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[4]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[12]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[12]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[20]\, Y
         => \MemorySynchronizer_0/N_1079\);
    
    \MemorySynchronizer_0/ConfigReg[15]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[15]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[12]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[1]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[12]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[12]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_23\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[16]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[16]\);
    
    \MemorySynchronizer_0/numberofnewavails_0_sqmuxa_0_a2_0_a2\ : 
        CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/APBState_Z[1]\, B => 
        \MemorySynchronizer_0/N_2567\, C => 
        \MemorySynchronizer_0/N_2586\, Y => 
        \MemorySynchronizer_0/numberofnewavails_0_sqmuxa\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[28]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[28]\);
    
    \STAMP_0/un85_paddr_3_RNIBFJK\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \STAMP_0/un85_paddr_3_Z\, B => 
        debug_led_net_0, C => \STAMP_0/component_state_Z[3]\, D
         => sb_sb_0_STAMP_PWRITE, Y => 
        \STAMP_0/un1_presetn_inv_i\);
    
    \STAMP_0/spi_request_for[1]\ : SLE
      port map(D => \STAMP_0/N_568_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_4_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_request_for_Z[1]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[1]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/N_2588\, B => 
        \MemorySynchronizer_0/N_2597\, C => 
        \MemorySynchronizer_0/TimeStampReg_Z[1]\, D => 
        \MemorySynchronizer_0/ConfigReg_Z[1]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[1]\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_1\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[1]\, 
        B => \MemorySynchronizer_0/un104_in_enable_0\, C => 
        \MemorySynchronizer_0/un104_in_enable_1\, D => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_Y\, 
        FCI => ADLIB_GND0, S => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[0]\, CC
         => NET_CC_CONFIG538, P => NET_CC_CONFIG536, UB => 
        NET_CC_CONFIG537);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[13]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_m_0_0[13]\, B
         => ENABLE_MEMORY_LED_c, C => \sb_sb_0_STAMP_PWDATA[13]\, 
        D => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, 
        Y => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[13]\);
    
    \STAMP_0/spi/count_cry[22]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[22]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[21]\, S => 
        \STAMP_0/spi/count_s[22]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[22]\, CC => NET_CC_CONFIG991, P
         => NET_CC_CONFIG989, UB => NET_CC_CONFIG990);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_i_i_a2_fast[0]\ : 
        CFG1
      generic map(INIT => "01")

      port map(A => \MemorySynchronizer_0/temp_1_cry_0_Y\, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_i_i_a2_fast_Z[0]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10[31]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \sb_sb_0_STAMP_PADDR[5]\, B => 
        \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[3]\, Y => 
        \MemorySynchronizer_0/N_2561\);
    
    \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_2_i\ : CFG3
      generic map(INIT => x"FD")

      port map(A => stamp0_ready_temp_c, B => 
        \STAMP_0/request_resync_0_sqmuxa\, C => 
        \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_1\, Y => 
        \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_2_i_Z\);
    
    \STAMP_0/spi/clk_toggles_lm_0[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/spi/ss_n_buffer_1_sqmuxa\, B => 
        \STAMP_0/spi/clk_toggles_s[1]\, Y => 
        \STAMP_0/spi/clk_toggles_lm[1]\);
    
    \STAMP_0/measurement_temp[11]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[27]\);
    
    \STAMP_0/component_state[0]\ : SLE
      port map(D => \STAMP_0/N_487_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/component_state_Z[0]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_10\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[10]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_9_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[22]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_10_Z\, CC
         => NET_CC_CONFIG327, P => NET_CC_CONFIG325, UB => 
        NET_CC_CONFIG326);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_18\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[18]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[18]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_17\, S => 
        \MemorySynchronizer_0/temp_1[18]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_18\, CC => 
        NET_CC_CONFIG253, P => NET_CC_CONFIG251, UB => 
        NET_CC_CONFIG252);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_1\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/CLK1_net\, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/PENABLE_net\, IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[17]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_17\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[8]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[8]\, B => 
        \sb_sb_0_STAMP_PWDATA[8]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[8]\);
    
    AFLSDF_INV_95 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_34\, Y => 
        \AFLSDF_INV_95\);
    
    \STAMP_0/spi/state_RNI1POH1[0]\ : CFG4
      generic map(INIT => x"E200")

      port map(A => \STAMP_0/enable\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, D => debug_led_net_0, Y => 
        \STAMP_0/spi/N_37_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_50\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_54_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[12]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_54\);
    
    \STAMP_0/un1_pwdata[10]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[10]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => 
        \STAMP_0/un1_pwdata_Z[10]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[4]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_4\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[20]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_20_S\, 
        Y => \MemorySynchronizer_0/N_1513\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[30]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \MemorySynchronizer_0/N_2588\, B => 
        \MemorySynchronizer_0/N_2597\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[30]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[30]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[30]\);
    
    \STAMP_0/delay_counter_cry[12]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[12]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[11]\, S
         => \STAMP_0/delay_counter_s[12]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[12]\, CC => NET_CC_CONFIG431, 
        P => NET_CC_CONFIG429, UB => NET_CC_CONFIG430);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[18]\ : SLE
      port map(D => \STAMP_0_data_frame[50]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[18]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[26]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[26]\, B => 
        \MemorySynchronizer_0/un104_in_enable_26\, C => 
        \MemorySynchronizer_0/N_2574\, D => 
        \MemorySynchronizer_0/N_2577\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[26]\);
    
    \STAMP_0/spi/count[10]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[10]\);
    
    \MemorySynchronizer_0/waitingtimercounter[14]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[14]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_52_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[14]\);
    
    \STAMP_0/measurement_dms2_1_sqmuxa_0_a3\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \STAMP_0/apb_spi_finished_0_sqmuxa_1\, B => 
        debug_led_net_0, C => \STAMP_0/spi_request_for_Z[1]\, D
         => \STAMP_0/spi_request_for_Z[0]\, Y => 
        \STAMP_0/measurement_dms2_1_sqmuxa\);
    
    \STAMP_0/delay_counter_lm_0[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[26]\, Y => 
        \STAMP_0/delay_counter_lm[26]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_70\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4]\, 
        IPC => OPEN);
    
    \STAMP_0/status_async_cycles[3]\ : SLE
      port map(D => \STAMP_0/status_async_cycles_lm[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/status_async_cycles_1_sqmuxa_1_i_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[6]\);
    
    \STAMP_0/delay_counter_lm_0[18]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[18]\, Y => 
        \STAMP_0/delay_counter_lm[18]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_10[20]\ : 
        CFG2
      generic map(INIT => x"1")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[0]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[5]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_10_Z[20]\);
    
    \STAMP_0/un1_spi_rx_data_0[23]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[23]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[23]\, Y
         => \STAMP_0/N_606\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_21\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[21]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_20_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[11]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_21_Z\, CC
         => NET_CC_CONFIG360, P => NET_CC_CONFIG358, UB => 
        NET_CC_CONFIG359);
    
    \MemorySynchronizer_0/un1_nreset_20_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_47\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_20_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_20_rs_Z\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[26]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB0_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[26]\);
    
    \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_3_i_0_a2_1\ : 
        CFG4
      generic map(INIT => x"4000")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[3]\, D => \sb_sb_0_STAMP_PADDR[5]\, 
        Y => \MemorySynchronizer_0/N_2586\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[24]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[24]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[24]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[24]\);
    
    AFLSDF_INV_29 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_29\);
    
    ResetAND : CFG2
      generic map(INIT => x"8")

      port map(A => sb_sb_0_POWER_ON_RESET_N, B => 
        sb_sb_0_GPIO_4_M2F, Y => NN_1);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2\ : 
        CFG4
      generic map(INIT => x"AE00")

      port map(A => STAMP_0_new_avail, B => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_28_Z\, 
        C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2_1\, 
        D => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, Y
         => \MemorySynchronizer_0/N_140_2\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[31]\ : SLE
      port map(D => \STAMP_0_data_frame[63]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[31]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[17]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[17]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[17]\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[17]\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[17]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[1]\ : SLE
      port map(D => \STAMP_0_data_frame[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[1]\);
    
    \STAMP_0/spi/busy\ : SLE
      port map(D => \STAMP_0/spi/busy_7\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_busy\);
    
    AFLSDF_INV_89 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_47\, Y => 
        \AFLSDF_INV_89\);
    
    \STAMP_0/spi/tx_buffer_RNO[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[13]\, B => 
        \STAMP_0/spi/tx_buffer_Z[12]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_122\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[28]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[28]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[28]\);
    
    \STAMP_0/config[22]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[22]\);
    
    AFLSDF_INV_27 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_27\);
    
    \STAMP_0/spi/tx_buffer[7]\ : SLE
      port map(D => \STAMP_0/spi/N_128\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[7]\);
    
    \STAMP_0/spi_enable\ : SLE
      port map(D => \STAMP_0/spi_enable_RNO_Z\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/N_244\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/enable\);
    
    \MemorySynchronizer_0/waitingtimercounter[5]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_5_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[5]\);
    
    \MemorySynchronizer_0/un1_nreset_32\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[2]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_32_i\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_CC_0\ : 
        CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => CI_TO_CO100, P(0) => 
        ADLIB_GND0, P(1) => NET_CC_CONFIG102, P(2) => 
        NET_CC_CONFIG105, P(3) => NET_CC_CONFIG108, P(4) => 
        NET_CC_CONFIG111, P(5) => NET_CC_CONFIG114, P(6) => 
        NET_CC_CONFIG117, P(7) => NET_CC_CONFIG120, P(8) => 
        NET_CC_CONFIG123, P(9) => NET_CC_CONFIG126, P(10) => 
        NET_CC_CONFIG129, P(11) => NET_CC_CONFIG132, UB(0) => 
        ADLIB_VCC1, UB(1) => NET_CC_CONFIG103, UB(2) => 
        NET_CC_CONFIG106, UB(3) => NET_CC_CONFIG109, UB(4) => 
        NET_CC_CONFIG112, UB(5) => NET_CC_CONFIG115, UB(6) => 
        NET_CC_CONFIG118, UB(7) => NET_CC_CONFIG121, UB(8) => 
        NET_CC_CONFIG124, UB(9) => NET_CC_CONFIG127, UB(10) => 
        NET_CC_CONFIG130, UB(11) => NET_CC_CONFIG133, CC(0) => 
        nc252, CC(1) => NET_CC_CONFIG104, CC(2) => 
        NET_CC_CONFIG107, CC(3) => NET_CC_CONFIG110, CC(4) => 
        NET_CC_CONFIG113, CC(5) => NET_CC_CONFIG116, CC(6) => 
        NET_CC_CONFIG119, CC(7) => NET_CC_CONFIG122, CC(8) => 
        NET_CC_CONFIG125, CC(9) => NET_CC_CONFIG128, CC(10) => 
        NET_CC_CONFIG131, CC(11) => NET_CC_CONFIG134);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_4\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_5\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_3_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[5]\, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_4_Z\, 
        CC => NET_CC_CONFIG1035, P => NET_CC_CONFIG1033, UB => 
        NET_CC_CONFIG1034);
    
    AFLSDF_INV_87 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_35\, Y => 
        \AFLSDF_INV_87\);
    
    \stamp0_ready_dms2_ibuf/U0/U_IOPAD\ : sdf_IOPAD_IN
      port map(PAD => stamp0_ready_dms2, Y => 
        \stamp0_ready_dms2_ibuf/U0/YIN1\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_239\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_23\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[23]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[23]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_22\, S => 
        \MemorySynchronizer_0/temp_1[23]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_23\, CC => 
        NET_CC_CONFIG268, P => NET_CC_CONFIG266, UB => 
        NET_CC_CONFIG267);
    
    \STAMP_0/spi/count[14]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[14]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_2\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[2]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[2]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_1_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_2_Z\, CC => 
        NET_CC_CONFIG829, P => NET_CC_CONFIG827, UB => 
        NET_CC_CONFIG828);
    
    \MemorySynchronizer_0/un1_nreset_8\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[29]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_8_i\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[26]\ : SLE
      port map(D => \STAMP_0_data_frame[58]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[26]\);
    
    \STAMP_0/spi/rx_buffer[1]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[1]\);
    
    \STAMP_0/delay_counter[0]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[0]\);
    
    \STAMP_0/new_avail\ : SLE
      port map(D => \STAMP_0/new_avail_0_sqmuxa_1\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_new_avail_1_sqmuxa_3_i_0_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => STAMP_0_new_avail);
    
    \STAMP_0/component_state_ns_0_i_o2_0[0]\ : CFG3
      generic map(INIT => x"FD")

      port map(A => \STAMP_0/component_state_Z[2]\, B => 
        sb_sb_0_STAMP_PENABLE, C => \STAMP_0/apb_is_atomic_Z\, Y
         => \STAMP_0/N_167\);
    
    \STAMP_0/spi/tx_buffer[0]\ : SLE
      port map(D => \STAMP_0/spi/N_333\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[0]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[20]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[20]\);
    
    \STAMP_0/async_prescaler_count[11]\ : SLE
      port map(D => \STAMP_0/async_prescaler_count_5_Z[11]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \STAMP_0/async_prescaler_count_Z[11]\);
    
    AFLSDF_INV_1 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_1\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_27\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[27]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_26_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_27_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_27_Z\, CC
         => NET_CC_CONFIG806, P => NET_CC_CONFIG804, UB => 
        NET_CC_CONFIG805);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[4]\ : SLE
      port map(D => \STAMP_0_data_frame[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[4]\);
    
    \MemorySynchronizer_0/un1_nreset_23_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_60_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_23_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_23_rs_Z\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[24]\ : SLE
      port map(D => \STAMP_0_data_frame[56]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[24]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_201\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[23]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[23]\, B => 
        \sb_sb_0_STAMP_PWDATA[23]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[23]\);
    
    AFLSDF_INV_58 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_58\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_9\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_10\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_8_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[10]\, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_9_Z\, 
        CC => NET_CC_CONFIG1050, P => NET_CC_CONFIG1048, UB => 
        NET_CC_CONFIG1049);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_30\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[30]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_29_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[2]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_FCNET1\, 
        CC => NET_CC_CONFIG387, P => NET_CC_CONFIG385, UB => 
        NET_CC_CONFIG386);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_19\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[19]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_18_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_19_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_19_Z\, CC
         => NET_CC_CONFIG782, P => NET_CC_CONFIG780, UB => 
        NET_CC_CONFIG781);
    
    \MemorySynchronizer_0/SynchStatusReg2_RNO[26]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \MemorySynchronizer_0/temp_1_cry_0_Y\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[26]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[26]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_30\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[30]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_29_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_30_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_30_Z\, 
        CC => NET_CC_CONFIG717, P => NET_CC_CONFIG715, UB => 
        NET_CC_CONFIG716);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_31[20]\ : 
        CFG4
      generic map(INIT => x"2000")

      port map(A => \MemorySynchronizer_0/un151_in_enable\, B => 
        \MemorySynchronizer_0/N_2328\, C => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_27_Z[20]\, 
        D => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_28_Z[20]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_31_Z[20]\);
    
    \STAMP_0/spi_tx_data[14]\ : SLE
      port map(D => \STAMP_0/N_267_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[14]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[8]\ : SLE
      port map(D => \STAMP_0_data_frame[40]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[8]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[20]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[20]\);
    
    \MMUART_0_RXD_F2M_ibuf/U0/U_IOINFF\ : IOINFF_BYPASS
      port map(A => \MMUART_0_RXD_F2M_ibuf/U0/YIN1\, Y => 
        \MMUART_0_RXD_F2M_ibuf/U0/YIN\);
    
    \STAMP_0/measurement_temp[5]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[21]\);
    
    \STAMP_0/delay_counter[16]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[16]\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_20\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[14]\, B => 
        \MemorySynchronizer_0/un120_in_enable_i_A[15]\, C => 
        \MemorySynchronizer_0/un120_in_enable_i_A[16]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[17]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_20_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[22]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_22_S\, 
        Y => \MemorySynchronizer_0/N_1501\);
    
    \STAMP_0/un1_spi_rx_data_1[22]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[54]\, B => 
        \STAMP_0/dummy_Z[22]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_639\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_19\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[10]\, B => 
        \MemorySynchronizer_0/un120_in_enable_i_A[11]\, C => 
        \MemorySynchronizer_0/un120_in_enable_i_A[12]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[13]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_19_Z\);
    
    
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_1_1_RNISF2T1[4]\ : 
        CFG4
      generic map(INIT => x"1300")

      port map(A => \MemorySynchronizer_0/N_140_2\, B => 
        \MemorySynchronizer_0/N_6\, C => 
        \MemorySynchronizer_0/N_2330\, D => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_1_1_Z[4]\, 
        Y => \MemorySynchronizer_0/N_2510\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[24]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[24]\, B => 
        \sb_sb_0_STAMP_PWDATA[24]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[24]\);
    
    \STAMP_0/apb_is_reset\ : SLE
      port map(D => \sb_sb_0_STAMP_PADDR[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/apb_is_atomic_0_sqmuxa\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/apb_is_reset_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_167\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg[3]\ : SLE
      port map(D => \MemorySynchronizer_0/SynchStatusReg_168[1]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, 
        EN => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[3]\);
    
    \MemorySynchronizer_0/SynchStatusReg[6]\ : SLE
      port map(D => \MemorySynchronizer_0/SynchStatusReg_168[4]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, 
        EN => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[6]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[3]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[3]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[3]\, D => 
        \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[3]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[20]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[20]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[20]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[20]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[20]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[20]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[16]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[16]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[16]\, C => 
        \MemorySynchronizer_0/N_2593\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[16]\);
    
    \STAMP_0/spi/tx_buffer[15]\ : SLE
      port map(D => \STAMP_0/spi/N_120\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[15]\);
    
    \MemorySynchronizer_0/TimeStampReg[0]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[0]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[0]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[2]\ : SLE
      port map(D => \STAMP_0_data_frame[34]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[2]\);
    
    \stamp0_spi_mosi_obuft/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \stamp0_spi_mosi_obuft/U0/DOUT1\, Y => 
        \stamp0_spi_mosi_obuft/U0/DOUT\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[29]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[29]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1062\, Y => 
        \MemorySynchronizer_0/N_1093\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_1[28]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[29]\, 
        B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_16_0_Z[28]\, C
         => \MemorySynchronizer_0/N_1182\, Y => 
        \MemorySynchronizer_0/N_1163\);
    
    \MemorySynchronizer_0/SynchStatusReg[28]\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg_152_e2\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[28]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_25\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[25]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_24_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[7]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_25_Z\, CC
         => NET_CC_CONFIG372, P => NET_CC_CONFIG370, UB => 
        NET_CC_CONFIG371);
    
    \STAMP_0/un1_spi_rx_data_0[8]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[8]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[8]\, Y
         => \STAMP_0/N_591\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[17]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[17]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[17]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_43\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net\, 
        IPC => OPEN);
    
    \STAMP_0/drdy_flank_detected_dms1_RNO\ : CFG1
      generic map(INIT => "01")

      port map(A => stamp0_ready_dms1_c, Y => 
        \STAMP_0/stamp0_ready_dms1_c_i\);
    
    \STAMP_0/component_state_ns_0_0_a3_1[2]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/apb_spi_finished_Z\, B => 
        \STAMP_0/component_state_Z[0]\, C => 
        \STAMP_0/component_state_Z[3]\, Y => 
        \STAMP_0/component_state_ns_0_0_a3_1_Z[2]\);
    
    \MISO_ibuf/U0/U_IOINFF\ : IOINFF_BYPASS
      port map(A => \MISO_ibuf/U0/YIN1\, Y => \MISO_ibuf/U0/YIN\);
    
    AFLSDF_INV_40 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_40\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_20_x\ : 
        CFG3
      generic map(INIT => x"01")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[14]\, B => 
        \MemorySynchronizer_0/un120_in_enable_i_A[15]\, C => 
        \MemorySynchronizer_0/un120_in_enable_i_A[16]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_20_x_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_a2_0[0]\ : 
        CFG2
      generic map(INIT => x"4")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, B => 
        \MemorySynchronizer_0/SynchStatusReg_Z[2]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_a2_0_Z[0]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[28]\ : SLE
      port map(D => \STAMP_0_data_frame[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[28]\);
    
    \MemorySynchronizer_0/MemorySyncState[4]\ : SLE
      port map(D => \MemorySynchronizer_0/MemorySyncState_ns[1]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, 
        EN => ENABLE_MEMORY_LED_c, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/MemorySyncState_Z[4]\);
    
    \STAMP_0/un5_async_prescaler_count_cry_7\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[7]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_6_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_7_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_7_Z\, CC
         => NET_CC_CONFIG501, P => NET_CC_CONFIG499, UB => 
        NET_CC_CONFIG500);
    
    \MemorySynchronizer_0/resettimercounter[3]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[3]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_31_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[3]\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_39\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[13]\, B => 
        \MemorySynchronizer_0/un104_in_enable_12\, C => 
        \MemorySynchronizer_0/un104_in_enable_13\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[12]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[5]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[6]\, CC
         => NET_CC_CONFIG556, P => NET_CC_CONFIG554, UB => 
        NET_CC_CONFIG555);
    
    \STAMP_0/un45_async_state_cry_2\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \STAMP_0/config_Z[26]\, B => 
        \STAMP_0_data_frame[5]\, C => ADLIB_GND0, D => ADLIB_GND0, 
        FCI => \STAMP_0/un45_async_state_cry_1_Z\, S => OPEN, Y
         => OPEN, FCO => \STAMP_0/un45_async_state_cry_2_Z\, CC
         => NET_CC_CONFIG522, P => NET_CC_CONFIG520, UB => 
        NET_CC_CONFIG521);
    
    \MemorySynchronizer_0/resynctimercounter[25]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1097\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[25]\);
    
    \STAMP_0/config[10]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[10]\);
    
    \STAMP_0/spi/count_cry[9]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[9]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[8]\, S => 
        \STAMP_0/spi/count_s[9]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[9]\, CC => NET_CC_CONFIG952, P
         => NET_CC_CONFIG950, UB => NET_CC_CONFIG951);
    
    \STAMP_0/un52_paddr_2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \sb_sb_0_STAMP_PADDR[9]\, B => 
        \sb_sb_0_STAMP_PADDR[7]\, C => \STAMP_0/un52_paddr_2_Z\, 
        D => \STAMP_0/un52_paddr_5_Z\, Y => 
        \STAMP_0/un52_paddr_2_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[9]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \MemorySynchronizer_0/N_2585\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[9]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[9]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[9]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_216\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[17]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[17]\);
    
    \STAMP_0/delay_counter[5]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[5]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[27]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[27]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[5]\, Y => 
        \MemorySynchronizer_0/N_1064\);
    
    \MemorySynchronizer_0/waitingtimercounter[17]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[17]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_24_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[17]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[24]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_24_S\, 
        Y => \MemorySynchronizer_0/N_2418\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[22]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[22]\);
    
    \MemorySynchronizer_0/un1_nreset_41_0_a3\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[12]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_41_i\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_31_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[19]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_31\);
    
    \STAMP_0/un1_spi_rx_data_0[20]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[20]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[20]\, Y
         => \STAMP_0/N_603\);
    
    \STAMP_0/spi/rx_buffer_0_sqmuxa_1_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \STAMP_0/spi/N_30\, B => 
        \STAMP_0/spi/ss_n_buffer_Z[0]\, C => debug_led_net_0, D
         => \STAMP_0/spi/N_63\, Y => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_22\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[22]\, B => 
        \MemorySynchronizer_0/un120_in_enable_i_A[23]\, C => 
        \MemorySynchronizer_0/un120_in_enable_i_A[24]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[25]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_22_Z\);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.un151_in_enablelto30_19\ : 
        CFG3
      generic map(INIT => x"FE")

      port map(A => \MemorySynchronizer_0/temp_1[29]\, B => 
        \MemorySynchronizer_0/temp_1[30]\, C => 
        \MemorySynchronizer_0/un151_in_enablelto30_13\, Y => 
        \MemorySynchronizer_0/un151_in_enablelto30_19\);
    
    \STAMP_0/un5_async_prescaler_count_cry_3\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[3]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_2_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_3_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_3_Z\, CC
         => NET_CC_CONFIG489, P => NET_CC_CONFIG487, UB => 
        NET_CC_CONFIG488);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.un151_in_enablelto31\ : 
        CFG4
      generic map(INIT => x"E0F0")

      port map(A => 
        \MemorySynchronizer_0/un151_in_enablelto30_19\, B => 
        \MemorySynchronizer_0/un151_in_enablelto30_23\, C => 
        \MemorySynchronizer_0/temp_1_cry_30\, D => 
        \MemorySynchronizer_0/un151_in_enablelto31_1\, Y => 
        \MemorySynchronizer_0/un151_in_enable\);
    
    \STAMP_0/un1_spi_rx_data_2[24]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_607\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, C => \STAMP_0/N_641\, Y
         => \STAMP_0/N_674\);
    
    \STAMP_0/delay_counter[8]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[8]\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_16\ : CFG4
      generic map(INIT => x"0010")

      port map(A => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_2_S\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_3_S\, 
        C => \MemorySynchronizer_0/resettimercounter_Z[0]\, D => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_1_S\, Y
         => \MemorySynchronizer_0/un6_in_enable_0_a3_16_Z\);
    
    \STAMP_0/config[23]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[23]\);
    
    \MMUART_0_TXD_M2F_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \MMUART_0_TXD_M2F_obuf/U0/DOUT1\, Y => 
        \MMUART_0_TXD_M2F_obuf/U0/DOUT\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[10]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[10]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[22]\, Y
         => \MemorySynchronizer_0/N_1081\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_212\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/MemorySyncState_ns_i_0_i[3]\ : CFG4
      generic map(INIT => x"A200")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => \MemorySynchronizer_0/N_2313\, C => 
        \MemorySynchronizer_0/un1_in_enable_2_0_0_a2_0_Z\, D => 
        \MemorySynchronizer_0/N_140_2\, Y => 
        \MemorySynchronizer_0/N_304\);
    
    AFLSDF_INV_91 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_91\);
    
    \MemorySynchronizer_0/ConfigReg[16]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[16]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_30\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[30]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_29_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_30_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_30_Z\, CC
         => NET_CC_CONFIG815, P => NET_CC_CONFIG813, UB => 
        NET_CC_CONFIG814);
    
    \MemorySynchronizer_0/SynchStatusReg[24]\ : SLE
      port map(D => \MemorySynchronizer_0/N_215_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[24]\);
    
    \MemorySynchronizer_0/APBState[1]\ : SLE
      port map(D => \MemorySynchronizer_0/APBState_ns[1]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/APBState_Z[1]\);
    
    \STAMP_0/delay_counter_cry[21]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[21]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[20]\, S
         => \STAMP_0/delay_counter_s[21]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[21]\, CC => NET_CC_CONFIG458, 
        P => NET_CC_CONFIG456, UB => NET_CC_CONFIG457);
    
    \STAMP_0/spi_tx_data_RNO[15]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[15]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_268_i\);
    
    \MemorySynchronizer_0/PRDATA[7]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[7]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[7]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[29]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[29]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[29]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_1\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => \sb_sb_0_STAMP_PADDR[4]\, B => 
        \sb_sb_0_STAMP_PADDR[2]\, Y => 
        \MemorySynchronizer_0/N_2567\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_8[28]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_2564\, C => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_2574\);
    
    \MemorySynchronizer_0/ResetTimerValueReg_RNINBVC[15]\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[15]\, B => 
        NN_1, Y => \MemorySynchronizer_0/N_1979_i\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[26]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[26]\, B => 
        \sb_sb_0_STAMP_PWDATA[26]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[26]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_0_CC_1\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO293, CO => CI_TO_CO294, P(0) => 
        NET_CC_CONFIG331, P(1) => NET_CC_CONFIG334, P(2) => 
        NET_CC_CONFIG337, P(3) => NET_CC_CONFIG340, P(4) => 
        NET_CC_CONFIG343, P(5) => NET_CC_CONFIG346, P(6) => 
        NET_CC_CONFIG349, P(7) => NET_CC_CONFIG352, P(8) => 
        NET_CC_CONFIG355, P(9) => NET_CC_CONFIG358, P(10) => 
        NET_CC_CONFIG361, P(11) => NET_CC_CONFIG364, UB(0) => 
        NET_CC_CONFIG332, UB(1) => NET_CC_CONFIG335, UB(2) => 
        NET_CC_CONFIG338, UB(3) => NET_CC_CONFIG341, UB(4) => 
        NET_CC_CONFIG344, UB(5) => NET_CC_CONFIG347, UB(6) => 
        NET_CC_CONFIG350, UB(7) => NET_CC_CONFIG353, UB(8) => 
        NET_CC_CONFIG356, UB(9) => NET_CC_CONFIG359, UB(10) => 
        NET_CC_CONFIG362, UB(11) => NET_CC_CONFIG365, CC(0) => 
        NET_CC_CONFIG333, CC(1) => NET_CC_CONFIG336, CC(2) => 
        NET_CC_CONFIG339, CC(3) => NET_CC_CONFIG342, CC(4) => 
        NET_CC_CONFIG345, CC(5) => NET_CC_CONFIG348, CC(6) => 
        NET_CC_CONFIG351, CC(7) => NET_CC_CONFIG354, CC(8) => 
        NET_CC_CONFIG357, CC(9) => NET_CC_CONFIG360, CC(10) => 
        NET_CC_CONFIG363, CC(11) => NET_CC_CONFIG366);
    
    AFLSDF_INV_69 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_51\, Y => 
        \AFLSDF_INV_69\);
    
    \stamp0_spi_temp_cs_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \stamp0_spi_temp_cs_obuf/U0/EOUT1\, Y => 
        \stamp0_spi_temp_cs_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/waitingtimercounter[20]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[20]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_62_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[20]\);
    
    AFLSDF_INV_67 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_67\);
    
    \MemorySynchronizer_0/ConfigReg[2]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[2]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[4]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[4]\);
    
    \MemorySynchronizer_0/MemorySyncState[0]\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/MemorySyncStatece_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/MemorySyncState_Z[0]\);
    
    \STAMP_0/un1_spi_rx_data_0[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[5]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[5]\, Y
         => \STAMP_0/N_588\);
    
    \STAMP_0/un1_presetn_inv_4_i_0\ : CFG3
      generic map(INIT => x"C4")

      port map(A => \STAMP_0/N_219\, B => debug_led_net_0, C => 
        \STAMP_0/N_361\, Y => \STAMP_0/un1_presetn_inv_4_i_0_Z\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_7\ : CFG4
      generic map(INIT => x"0035")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_Z[2]\, B => 
        \MemorySynchronizer_0/resynctimercounter_1[30]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, D
         => \MemorySynchronizer_0/N_1076\, Y => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_7_Z\);
    
    \STAMP_0/spi/clk_toggles_lm_0[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/spi/ss_n_buffer_1_sqmuxa\, B => 
        \STAMP_0/spi/clk_toggles_s[3]\, Y => 
        \STAMP_0/spi/clk_toggles_lm[3]\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2_N_2L1\ : 
        CFG4
      generic map(INIT => x"BFFF")

      port map(A => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2_N_2L1_1_Z\, 
        B => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[15]\, C
         => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_22_Z\, 
        D => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_23_Z\, 
        Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2_1\);
    
    \MemorySynchronizer_0/un1_nreset_27\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[27]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_27_i\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[8]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[8]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[8]\, C => 
        \MemorySynchronizer_0/N_2593\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[8]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_44_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_55\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_44_set_Z\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[19]\ : SLE
      port map(D => \STAMP_0_data_frame[51]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[19]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[21]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[21]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[21]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[21]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_3\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[18]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[18]\);
    
    \STAMP_0/un1_spi_rx_data_i_m2_0[30]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame[30]\, B => 
        \STAMP_0/config_Z[30]\, C => \sb_sb_0_STAMP_PADDR[8]\, Y
         => \STAMP_0/N_218\);
    
    \stamp0_spi_temp_cs_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \stamp0_spi_temp_cs_obuf/U0/DOUT1\, Y => 
        \stamp0_spi_temp_cs_obuf/U0/DOUT\);
    
    \STAMP_0/PRDATA[25]\ : SLE
      port map(D => \STAMP_0/N_675\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_56\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[25]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[9]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[9]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1082\, Y => 
        \MemorySynchronizer_0/N_1113\);
    
    \MemorySynchronizer_0/resettimercounter[27]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_27_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[27]\);
    
    \STAMP_0/status_dms2_overwrittenVal\ : SLE
      port map(D => \STAMP_0/N_117_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_new_avail_0_sqmuxa_3_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[11]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[19]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[19]\, B => 
        \sb_sb_0_STAMP_PWDATA[19]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[19]\);
    
    \MemorySynchronizer_0/resynctimercounter[5]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1117\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[5]\);
    
    \MemorySynchronizer_0/N_21_i_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_57\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_21_i_set_Z\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_42_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[30]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_42\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[18]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[18]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[17]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[18]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[18]\, CC
         => NET_CC_CONFIG60, P => NET_CC_CONFIG58, UB => 
        NET_CC_CONFIG59);
    
    \MemorySynchronizer_0/ConfigReg[20]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[20]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_20\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[20]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_19_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_20_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_20_Z\, CC
         => NET_CC_CONFIG785, P => NET_CC_CONFIG783, UB => 
        NET_CC_CONFIG784);
    
    \MemorySynchronizer_0/un1_nreset_48_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_46_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_48_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_48_rs_Z\);
    
    \STAMP_0/spi_tx_data[9]\ : SLE
      port map(D => \STAMP_0/N_289_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[9]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_51\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[5]\ : SLE
      port map(D => \STAMP_0_data_frame[37]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[5]\);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_23\ : 
        CFG4
      generic map(INIT => x"1000")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[7]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[9]\, C => 
        STAMP_0_new_avail, D => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_2_Z[20]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_23_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_0[20]\ : CFG2
      generic map(INIT => x"B")

      port map(A => 
        \MemorySynchronizer_0/un1_enabletimestampgen2_2_sn\, B
         => STAMP_0_new_avail, Y => \MemorySynchronizer_0/N_2328\);
    
    \STAMP_0/spi/count_lm_0[14]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[14]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[14]\);
    
    \MemorySynchronizer_0/un1_nreset_58_rs_RNI8PCH\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_2532_set_Z\, B => 
        \MemorySynchronizer_0/waitingtimercounterrs[8]\, C => 
        \MemorySynchronizer_0/un1_nreset_58_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[8]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[19]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[19]\, B => 
        \sb_sb_0_Memory_PRDATA[19]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[19]\);
    
    \STAMP_0/config[1]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[1]\);
    
    \MemorySynchronizer_0/resynctimercounter[17]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1105\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[17]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_71\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_4[3]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_3_S\, 
        Y => \MemorySynchronizer_0/N_1209\);
    
    \STAMP_0/spi_tx_data_RNO[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[5]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_293_i\);
    
    \MMUART_0_RXD_F2M_ibuf/U0/U_IOPAD\ : sdf_IOPAD_IN
      port map(PAD => MMUART_0_RXD_F2M, Y => 
        \MMUART_0_RXD_F2M_ibuf/U0/YIN1\);
    
    \STAMP_0/status_async_cycles_s_388\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0_data_frame[3]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => ADLIB_VCC1, S => 
        OPEN, Y => OPEN, FCO => 
        \STAMP_0/status_async_cycles_s_388_FCO\, CC => 
        NET_CC_CONFIG589, P => NET_CC_CONFIG587, UB => 
        NET_CC_CONFIG588);
    
    \MemorySynchronizer_0/PRDATA[19]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[19]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[19]\);
    
    AFLSDF_INV_4 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_4\);
    
    
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa_0_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/N_2567\, B => 
        \MemorySynchronizer_0/N_2586\, C => 
        \MemorySynchronizer_0/APBState_Z[1]\, D => 
        \sb_sb_0_STAMP_PWDATA[30]\, Y => 
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa\);
    
    \STAMP_0/config[15]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[15]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[27]\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \MemorySynchronizer_0/N_2577\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[27]\, C => 
        \MemorySynchronizer_0/un104_in_enable_27\, D => 
        \MemorySynchronizer_0/N_1411\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[27]\);
    
    \MemorySynchronizer_0/PRDATA[13]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[13]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa\ : CFG4
      generic map(INIT => x"0004")

      port map(A => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS[0]\, B => 
        sb_sb_0_STAMP_PSELx, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS_Z[2]\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS[1]\, Y => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_133\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15]\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/status_async_cycles_1_sqmuxa\ : CFG3
      generic map(INIT => x"02")

      port map(A => \STAMP_0/async_state_Z[0]\, B => 
        \STAMP_0/async_state_Z[1]\, C => 
        \STAMP_0/un1_async_prescaler_count\, Y => 
        \STAMP_0/status_async_cycles_1_sqmuxa_Z\);
    
    \STAMP_0/component_state[5]\ : SLE
      port map(D => \STAMP_0/N_100_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/component_state_Z[5]\);
    
    \RXSM_LO_ibuf/U0/U_IOINFF\ : IOINFF_BYPASS
      port map(A => \RXSM_LO_ibuf/U0/YIN1\, Y => 
        \RXSM_LO_ibuf/U0/YIN\);
    
    \STAMP_0/dummy[25]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_58\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[25]\);
    
    \STAMP_0/PRDATA[7]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[7]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[2]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[2]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[4]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[2]\);
    
    \STAMP_0/un1_component_state_13_i_o2\ : CFG2
      generic map(INIT => x"D")

      port map(A => \STAMP_0/N_111_i\, B => 
        \STAMP_0/config_Z[31]\, Y => \STAMP_0/N_164\);
    
    \STAMP_0/spi/count_cry[17]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[17]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[16]\, S => 
        \STAMP_0/spi/count_s[17]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[17]\, CC => NET_CC_CONFIG976, P
         => NET_CC_CONFIG974, UB => NET_CC_CONFIG975);
    
    \STAMP_0/spi/count[0]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[0]\);
    
    \STAMP_0/dummy_1_sqmuxa_4\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sb_sb_0_STAMP_PADDR[7]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/un52_paddr_2_0_Z\, 
        Y => \STAMP_0/dummy_1_sqmuxa_4_Z\);
    
    \MemorySynchronizer_0/un1_nreset_2_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_48\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_2_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_2_rs_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/INST_MSS_010_IP\ : 
        MSS_010_IP

              generic map(INIT => "00" & x"000000000000030000000000000000000000C00000000000000000000000000000000000000000000000000000000000C030000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFF82FAF09007C33C804000006092C0000003FFFFE4000000000024100000000F0F01C000001825F04010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem",
         RTC_MAIN_XTL_FREQ => 0.000000, RTC_MAIN_XTL_MODE => "",
         DDR_CLK_FREQ => 100.000000)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => sb_sb_0_GPIO_3_M2F, 
        CAN_TX_EBL_MGPIO4A_H2F_A => OPEN, 
        CAN_TX_EBL_MGPIO4A_H2F_B => sb_sb_0_GPIO_4_M2F, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => OPEN, COMMS_INT => OPEN, 
        CONFIG_PRESET_N => OPEN, EDAC_ERROR(7) => nc171, 
        EDAC_ERROR(6) => nc54, EDAC_ERROR(5) => nc286, 
        EDAC_ERROR(4) => nc307, EDAC_ERROR(3) => nc135, 
        EDAC_ERROR(2) => nc41, EDAC_ERROR(1) => nc100, 
        EDAC_ERROR(0) => nc404, F_FM0_RDATA(31) => nc270, 
        F_FM0_RDATA(30) => nc339, F_FM0_RDATA(29) => nc52, 
        F_FM0_RDATA(28) => nc251, F_FM0_RDATA(27) => nc186, 
        F_FM0_RDATA(26) => nc29, F_FM0_RDATA(25) => nc269, 
        F_FM0_RDATA(24) => nc118, F_FM0_RDATA(23) => nc412, 
        F_FM0_RDATA(22) => nc60, F_FM0_RDATA(21) => nc141, 
        F_FM0_RDATA(20) => nc311, F_FM0_RDATA(19) => nc276, 
        F_FM0_RDATA(18) => nc193, F_FM0_RDATA(17) => nc214, 
        F_FM0_RDATA(16) => nc298, F_FM0_RDATA(15) => nc282, 
        F_FM0_RDATA(14) => nc240, F_FM0_RDATA(13) => nc45, 
        F_FM0_RDATA(12) => nc53, F_FM0_RDATA(11) => nc121, 
        F_FM0_RDATA(10) => nc176, F_FM0_RDATA(9) => nc419, 
        F_FM0_RDATA(8) => nc360, F_FM0_RDATA(7) => nc220, 
        F_FM0_RDATA(6) => nc158, F_FM0_RDATA(5) => nc281, 
        F_FM0_RDATA(4) => nc209, F_FM0_RDATA(3) => nc427, 
        F_FM0_RDATA(2) => nc246, F_FM0_RDATA(1) => nc368, 
        F_FM0_RDATA(0) => nc351, F_FM0_READYOUT => OPEN, 
        F_FM0_RESP => OPEN, F_HM0_ADDR(31) => nc162, 
        F_HM0_ADDR(30) => nc11, F_HM0_ADDR(29) => nc272, 
        F_HM0_ADDR(28) => nc131, F_HM0_ADDR(27) => nc364, 
        F_HM0_ADDR(26) => nc254, F_HM0_ADDR(25) => nc267, 
        F_HM0_ADDR(24) => nc96, F_HM0_ADDR(23) => nc79, 
        F_HM0_ADDR(22) => nc441, F_HM0_ADDR(21) => nc226, 
        F_HM0_ADDR(20) => nc146, F_HM0_ADDR(19) => nc230, 
        F_HM0_ADDR(18) => nc89, F_HM0_ADDR(17) => nc119, 
        F_HM0_ADDR(16) => nc48, F_HM0_ADDR(15) => 
        \sb_sb_0/STAMP_PADDRS[15]\, F_HM0_ADDR(14) => 
        \sb_sb_0/STAMP_PADDRS[14]\, F_HM0_ADDR(13) => 
        \sb_sb_0/STAMP_PADDRS[13]\, F_HM0_ADDR(12) => 
        \sb_sb_0/STAMP_PADDRS[12]\, F_HM0_ADDR(11) => 
        \sb_sb_0_STAMP_PADDR[11]\, F_HM0_ADDR(10) => 
        \sb_sb_0_STAMP_PADDR[10]\, F_HM0_ADDR(9) => 
        \sb_sb_0_STAMP_PADDR[9]\, F_HM0_ADDR(8) => 
        \sb_sb_0_STAMP_PADDR[8]\, F_HM0_ADDR(7) => 
        \sb_sb_0_STAMP_PADDR[7]\, F_HM0_ADDR(6) => 
        \sb_sb_0_STAMP_PADDR[6]\, F_HM0_ADDR(5) => 
        \sb_sb_0_STAMP_PADDR[5]\, F_HM0_ADDR(4) => 
        \sb_sb_0_STAMP_PADDR[4]\, F_HM0_ADDR(3) => 
        \sb_sb_0_STAMP_PADDR[3]\, F_HM0_ADDR(2) => 
        \sb_sb_0_STAMP_PADDR[2]\, F_HM0_ADDR(1) => 
        \sb_sb_0_STAMP_PADDR[1]\, F_HM0_ADDR(0) => 
        \sb_sb_0_STAMP_PADDR[0]\, F_HM0_ENABLE => 
        sb_sb_0_STAMP_PENABLE, F_HM0_SEL => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx\, 
        F_HM0_SIZE(1) => nc437, F_HM0_SIZE(0) => nc271, 
        F_HM0_TRANS1 => OPEN, F_HM0_WDATA(31) => 
        \sb_sb_0_STAMP_PWDATA[31]\, F_HM0_WDATA(30) => 
        \sb_sb_0_STAMP_PWDATA[30]\, F_HM0_WDATA(29) => 
        \sb_sb_0_STAMP_PWDATA[29]\, F_HM0_WDATA(28) => 
        \sb_sb_0_STAMP_PWDATA[28]\, F_HM0_WDATA(27) => 
        \sb_sb_0_STAMP_PWDATA[27]\, F_HM0_WDATA(26) => 
        \sb_sb_0_STAMP_PWDATA[26]\, F_HM0_WDATA(25) => 
        \sb_sb_0_STAMP_PWDATA[25]\, F_HM0_WDATA(24) => 
        \sb_sb_0_STAMP_PWDATA[24]\, F_HM0_WDATA(23) => 
        \sb_sb_0_STAMP_PWDATA[23]\, F_HM0_WDATA(22) => 
        \sb_sb_0_STAMP_PWDATA[22]\, F_HM0_WDATA(21) => 
        \sb_sb_0_STAMP_PWDATA[21]\, F_HM0_WDATA(20) => 
        \sb_sb_0_STAMP_PWDATA[20]\, F_HM0_WDATA(19) => 
        \sb_sb_0_STAMP_PWDATA[19]\, F_HM0_WDATA(18) => 
        \sb_sb_0_STAMP_PWDATA[18]\, F_HM0_WDATA(17) => 
        \sb_sb_0_STAMP_PWDATA[17]\, F_HM0_WDATA(16) => 
        \sb_sb_0_STAMP_PWDATA[16]\, F_HM0_WDATA(15) => 
        \sb_sb_0_STAMP_PWDATA[15]\, F_HM0_WDATA(14) => 
        \sb_sb_0_STAMP_PWDATA[14]\, F_HM0_WDATA(13) => 
        \sb_sb_0_STAMP_PWDATA[13]\, F_HM0_WDATA(12) => 
        \sb_sb_0_STAMP_PWDATA[12]\, F_HM0_WDATA(11) => 
        \sb_sb_0_STAMP_PWDATA[11]\, F_HM0_WDATA(10) => 
        \sb_sb_0_STAMP_PWDATA[10]\, F_HM0_WDATA(9) => 
        \sb_sb_0_STAMP_PWDATA[9]\, F_HM0_WDATA(8) => 
        \sb_sb_0_STAMP_PWDATA[8]\, F_HM0_WDATA(7) => 
        \sb_sb_0_STAMP_PWDATA[7]\, F_HM0_WDATA(6) => 
        \sb_sb_0_STAMP_PWDATA[6]\, F_HM0_WDATA(5) => 
        \sb_sb_0_STAMP_PWDATA[5]\, F_HM0_WDATA(4) => 
        \sb_sb_0_STAMP_PWDATA[4]\, F_HM0_WDATA(3) => 
        \sb_sb_0_STAMP_PWDATA[3]\, F_HM0_WDATA(2) => 
        \sb_sb_0_STAMP_PWDATA[2]\, F_HM0_WDATA(1) => 
        \sb_sb_0_STAMP_PWDATA[1]\, F_HM0_WDATA(0) => 
        \sb_sb_0_STAMP_PWDATA[0]\, F_HM0_WRITE => 
        sb_sb_0_STAMP_PWRITE, FAB_CHRGVBUS => OPEN, 
        FAB_DISCHRGVBUS => OPEN, FAB_DMPULLDOWN => OPEN, 
        FAB_DPPULLDOWN => OPEN, FAB_DRVVBUS => OPEN, FAB_IDPULLUP
         => OPEN, FAB_OPMODE(1) => nc213, FAB_OPMODE(0) => nc421, 
        FAB_SUSPENDM => OPEN, FAB_TERMSEL => OPEN, FAB_TXVALID
         => OPEN, FAB_VCONTROL(3) => nc366, FAB_VCONTROL(2) => 
        nc300, FAB_VCONTROL(1) => nc126, FAB_VCONTROL(0) => nc195, 
        FAB_VCONTROLLOADM => OPEN, FAB_XCVRSEL(1) => nc188, 
        FAB_XCVRSEL(0) => nc242, FAB_XDATAOUT(7) => nc15, 
        FAB_XDATAOUT(6) => nc399, FAB_XDATAOUT(5) => nc308, 
        FAB_XDATAOUT(4) => nc236, FAB_XDATAOUT(3) => nc102, 
        FAB_XDATAOUT(2) => nc381, FAB_XDATAOUT(1) => nc304, 
        FAB_XDATAOUT(0) => nc3, FACC_GLMUX_SEL => OPEN, 
        FIC32_0_MASTER(1) => nc207, FIC32_0_MASTER(0) => nc47, 
        FIC32_1_MASTER(1) => nc90, FIC32_1_MASTER(0) => nc284, 
        FPGA_RESET_N => OPEN, GTX_CLK => OPEN, H2F_INTERRUPT(15)
         => nc222, H2F_INTERRUPT(14) => nc159, H2F_INTERRUPT(13)
         => nc431, H2F_INTERRUPT(12) => nc136, H2F_INTERRUPT(11)
         => nc241, H2F_INTERRUPT(10) => nc253, H2F_INTERRUPT(9)
         => nc178, H2F_INTERRUPT(8) => nc306, H2F_INTERRUPT(7)
         => nc215, H2F_INTERRUPT(6) => nc59, H2F_INTERRUPT(5) => 
        nc362, H2F_INTERRUPT(4) => nc221, H2F_INTERRUPT(3) => 
        nc371, H2F_INTERRUPT(2) => nc232, H2F_INTERRUPT(1) => 
        nc274, H2F_INTERRUPT(0) => nc18, H2F_NMI => OPEN, 
        H2FCALIB => OPEN, I2C0_SCL_MGPIO31B_H2F_A => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_B => LED_HEARTBEAT_c, 
        I2C0_SDA_MGPIO30B_H2F_A => OPEN, I2C0_SDA_MGPIO30B_H2F_B
         => LED_RECORDING_c, I2C1_SCL_MGPIO1A_H2F_A => OPEN, 
        I2C1_SCL_MGPIO1A_H2F_B => OPEN, I2C1_SDA_MGPIO0A_H2F_A
         => OPEN, I2C1_SDA_MGPIO0A_H2F_B => OPEN, MDCF => OPEN, 
        MDOENF => OPEN, MDOF => OPEN, MMUART0_CTS_MGPIO19B_H2F_A
         => OPEN, MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => nCS2_c, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => ENABLE_MEMORY_LED_c, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => nCS1_c, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => MMUART_0_TXD_M2F_c, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => OPEN, MPLL_LOCK => OPEN, 
        PER2_FABRIC_PADDR(15) => nc44, PER2_FABRIC_PADDR(14) => 
        nc117, PER2_FABRIC_PADDR(13) => nc418, 
        PER2_FABRIC_PADDR(12) => nc189, PER2_FABRIC_PADDR(11) => 
        nc164, PER2_FABRIC_PADDR(10) => nc148, 
        PER2_FABRIC_PADDR(9) => nc42, PER2_FABRIC_PADDR(8) => 
        nc231, PER2_FABRIC_PADDR(7) => nc191, 
        PER2_FABRIC_PADDR(6) => nc255, PER2_FABRIC_PADDR(5) => 
        nc442, PER2_FABRIC_PADDR(4) => nc283, 
        PER2_FABRIC_PADDR(3) => nc363, PER2_FABRIC_PADDR(2) => 
        nc341, PER2_FABRIC_PENABLE => OPEN, PER2_FABRIC_PSEL => 
        OPEN, PER2_FABRIC_PWDATA(31) => nc317, 
        PER2_FABRIC_PWDATA(30) => nc290, PER2_FABRIC_PWDATA(29)
         => nc17, PER2_FABRIC_PWDATA(28) => nc2, 
        PER2_FABRIC_PWDATA(27) => nc406, PER2_FABRIC_PWDATA(26)
         => nc302, PER2_FABRIC_PWDATA(25) => nc110, 
        PER2_FABRIC_PWDATA(24) => nc128, PER2_FABRIC_PWDATA(23)
         => nc414, PER2_FABRIC_PWDATA(22) => nc244, 
        PER2_FABRIC_PWDATA(21) => nc422, PER2_FABRIC_PWDATA(20)
         => nc321, PER2_FABRIC_PWDATA(19) => nc43, 
        PER2_FABRIC_PWDATA(18) => nc179, PER2_FABRIC_PWDATA(17)
         => nc157, PER2_FABRIC_PWDATA(16) => nc36, 
        PER2_FABRIC_PWDATA(15) => nc224, PER2_FABRIC_PWDATA(14)
         => nc296, PER2_FABRIC_PWDATA(13) => nc273, 
        PER2_FABRIC_PWDATA(12) => nc61, PER2_FABRIC_PWDATA(11)
         => nc104, PER2_FABRIC_PWDATA(10) => nc138, 
        PER2_FABRIC_PWDATA(9) => nc14, PER2_FABRIC_PWDATA(8) => 
        nc432, PER2_FABRIC_PWDATA(7) => nc357, 
        PER2_FABRIC_PWDATA(6) => nc285, PER2_FABRIC_PWDATA(5) => 
        nc429, PER2_FABRIC_PWDATA(4) => nc405, 
        PER2_FABRIC_PWDATA(3) => nc303, PER2_FABRIC_PWDATA(2) => 
        nc150, PER2_FABRIC_PWDATA(1) => nc365, 
        PER2_FABRIC_PWDATA(0) => nc331, PER2_FABRIC_PWRITE => 
        OPEN, RTC_MATCH => OPEN, SLEEPDEEP => OPEN, SLEEPHOLDACK
         => OPEN, SLEEPING => OPEN, SMBALERT_NO0 => OPEN, 
        SMBALERT_NO1 => OPEN, SMBSUS_NO0 => OPEN, SMBSUS_NO1 => 
        OPEN, SPI0_CLK_OUT => SCLK_c, SPI0_SDI_MGPIO5A_H2F_A => 
        OPEN, SPI0_SDI_MGPIO5A_H2F_B => OPEN, 
        SPI0_SDO_MGPIO6A_H2F_A => MOSI_c, SPI0_SDO_MGPIO6A_H2F_B
         => OPEN, SPI0_SS0_MGPIO7A_H2F_A => OPEN, 
        SPI0_SS0_MGPIO7A_H2F_B => OPEN, SPI0_SS1_MGPIO8A_H2F_A
         => OPEN, SPI0_SS1_MGPIO8A_H2F_B => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_A => OPEN, SPI0_SS2_MGPIO9A_H2F_B
         => OPEN, SPI0_SS3_MGPIO10A_H2F_A => OPEN, 
        SPI0_SS3_MGPIO10A_H2F_B => OPEN, SPI0_SS4_MGPIO19A_H2F_A
         => OPEN, SPI0_SS5_MGPIO20A_H2F_A => OPEN, 
        SPI0_SS6_MGPIO21A_H2F_A => OPEN, SPI0_SS7_MGPIO22A_H2F_A
         => OPEN, SPI1_CLK_OUT => OPEN, SPI1_SDI_MGPIO11A_H2F_A
         => OPEN, SPI1_SDI_MGPIO11A_H2F_B => OPEN, 
        SPI1_SDO_MGPIO12A_H2F_A => OPEN, SPI1_SDO_MGPIO12A_H2F_B
         => OPEN, SPI1_SS0_MGPIO13A_H2F_A => OPEN, 
        SPI1_SS0_MGPIO13A_H2F_B => OPEN, SPI1_SS1_MGPIO14A_H2F_A
         => OPEN, SPI1_SS1_MGPIO14A_H2F_B => OPEN, 
        SPI1_SS2_MGPIO15A_H2F_A => OPEN, SPI1_SS2_MGPIO15A_H2F_B
         => OPEN, SPI1_SS3_MGPIO16A_H2F_A => OPEN, 
        SPI1_SS3_MGPIO16A_H2F_B => OPEN, SPI1_SS4_MGPIO17A_H2F_A
         => OPEN, SPI1_SS5_MGPIO18A_H2F_A => OPEN, 
        SPI1_SS6_MGPIO23A_H2F_A => OPEN, SPI1_SS7_MGPIO24A_H2F_A
         => OPEN, TCGF(9) => nc196, TCGF(8) => nc234, TCGF(7) => 
        nc149, TCGF(6) => nc12, TCGF(5) => nc219, TCGF(4) => nc30, 
        TCGF(3) => nc243, TCGF(2) => nc187, TCGF(1) => nc65, 
        TCGF(0) => nc7, TRACECLK => OPEN, TRACEDATA(3) => nc292, 
        TRACEDATA(2) => nc439, TRACEDATA(1) => nc129, 
        TRACEDATA(0) => nc275, TX_CLK => OPEN, TX_ENF => OPEN, 
        TX_ERRF => OPEN, TXCTL_EN_RIF => OPEN, TXD_RIF(3) => nc8, 
        TXD_RIF(2) => nc223, TXD_RIF(1) => nc13, TXD_RIF(0) => 
        nc387, TXDF(7) => nc305, TXDF(6) => nc180, TXDF(5) => 
        nc26, TXDF(4) => nc291, TXDF(3) => nc177, TXDF(2) => 
        nc139, TXDF(1) => nc310, TXDF(0) => nc259, TXEV => OPEN, 
        WDOGTIMEOUT => OPEN, F_ARREADY_HREADYOUT1 => OPEN, 
        F_AWREADY_HREADYOUT0 => OPEN, F_BID(3) => nc403, F_BID(2)
         => nc245, F_BID(1) => nc233, F_BID(0) => nc163, 
        F_BRESP_HRESP0(1) => nc318, F_BRESP_HRESP0(0) => nc268, 
        F_BVALID => OPEN, F_RDATA_HRDATA01(63) => nc112, 
        F_RDATA_HRDATA01(62) => nc68, F_RDATA_HRDATA01(61) => 
        nc49, F_RDATA_HRDATA01(60) => nc377, F_RDATA_HRDATA01(59)
         => nc314, F_RDATA_HRDATA01(58) => nc217, 
        F_RDATA_HRDATA01(57) => nc170, F_RDATA_HRDATA01(56) => 
        nc91, F_RDATA_HRDATA01(55) => nc225, F_RDATA_HRDATA01(54)
         => nc5, F_RDATA_HRDATA01(53) => nc20, 
        F_RDATA_HRDATA01(52) => nc198, F_RDATA_HRDATA01(51) => 
        nc147, F_RDATA_HRDATA01(50) => nc350, 
        F_RDATA_HRDATA01(49) => nc316, F_RDATA_HRDATA01(48) => 
        nc391, F_RDATA_HRDATA01(47) => nc67, F_RDATA_HRDATA01(46)
         => nc289, F_RDATA_HRDATA01(45) => nc358, 
        F_RDATA_HRDATA01(44) => nc294, F_RDATA_HRDATA01(43) => 
        nc152, F_RDATA_HRDATA01(42) => nc127, 
        F_RDATA_HRDATA01(41) => nc103, F_RDATA_HRDATA01(40) => 
        nc428, F_RDATA_HRDATA01(39) => nc235, 
        F_RDATA_HRDATA01(38) => nc76, F_RDATA_HRDATA01(37) => 
        nc347, F_RDATA_HRDATA01(36) => nc208, 
        F_RDATA_HRDATA01(35) => nc354, F_RDATA_HRDATA01(34) => 
        nc140, F_RDATA_HRDATA01(33) => nc257, 
        F_RDATA_HRDATA01(32) => nc86, F_RDATA_HRDATA01(31) => 
        nc95, F_RDATA_HRDATA01(30) => nc327, F_RDATA_HRDATA01(29)
         => nc120, F_RDATA_HRDATA01(28) => nc424, 
        F_RDATA_HRDATA01(27) => nc165, F_RDATA_HRDATA01(26) => 
        nc356, F_RDATA_HRDATA01(25) => nc279, 
        F_RDATA_HRDATA01(24) => nc137, F_RDATA_HRDATA01(23) => 
        nc438, F_RDATA_HRDATA01(22) => nc64, F_RDATA_HRDATA01(21)
         => nc400, F_RDATA_HRDATA01(20) => nc19, 
        F_RDATA_HRDATA01(19) => nc380, F_RDATA_HRDATA01(18) => 
        nc369, F_RDATA_HRDATA01(17) => nc416, 
        F_RDATA_HRDATA01(16) => nc312, F_RDATA_HRDATA01(15) => 
        nc70, F_RDATA_HRDATA01(14) => nc388, F_RDATA_HRDATA01(13)
         => nc182, F_RDATA_HRDATA01(12) => nc62, 
        F_RDATA_HRDATA01(11) => nc337, F_RDATA_HRDATA01(10) => 
        nc199, F_RDATA_HRDATA01(9) => nc80, F_RDATA_HRDATA01(8)
         => nc130, F_RDATA_HRDATA01(7) => nc434, 
        F_RDATA_HRDATA01(6) => nc384, F_RDATA_HRDATA01(5) => 
        nc287, F_RDATA_HRDATA01(4) => nc98, F_RDATA_HRDATA01(3)
         => nc293, F_RDATA_HRDATA01(2) => nc249, 
        F_RDATA_HRDATA01(1) => nc114, F_RDATA_HRDATA01(0) => nc56, 
        F_RID(3) => nc370, F_RID(2) => nc105, F_RID(1) => nc386, 
        F_RID(0) => nc63, F_RLAST => OPEN, F_RRESP_HRESP1(1) => 
        nc415, F_RRESP_HRESP1(0) => nc352, F_RVALID => OPEN, 
        F_WREADY => OPEN, MDDR_FABRIC_PRDATA(15) => nc313, 
        MDDR_FABRIC_PRDATA(14) => nc309, MDDR_FABRIC_PRDATA(13)
         => nc378, MDDR_FABRIC_PRDATA(12) => nc172, 
        MDDR_FABRIC_PRDATA(11) => nc229, MDDR_FABRIC_PRDATA(10)
         => nc374, MDDR_FABRIC_PRDATA(9) => nc277, 
        MDDR_FABRIC_PRDATA(8) => nc97, MDDR_FABRIC_PRDATA(7) => 
        nc161, MDDR_FABRIC_PRDATA(6) => nc31, 
        MDDR_FABRIC_PRDATA(5) => nc340, MDDR_FABRIC_PRDATA(4) => 
        nc295, MDDR_FABRIC_PRDATA(3) => nc154, 
        MDDR_FABRIC_PRDATA(2) => nc376, MDDR_FABRIC_PRDATA(1) => 
        nc50, MDDR_FABRIC_PRDATA(0) => nc260, MDDR_FABRIC_PREADY
         => OPEN, MDDR_FABRIC_PSLVERR => OPEN, CAN_RXBUS_F2H_SCP
         => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net\, 
        CAN_TX_EBL_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net\, 
        CAN_TXBUS_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net\, 
        COLF => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/COLF_net\, 
        CRSF => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CRSF_net\, 
        F2_DMAREADY(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1]\, 
        F2_DMAREADY(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0]\, 
        F2H_INTERRUPT(15) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15]\, 
        F2H_INTERRUPT(14) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14]\, 
        F2H_INTERRUPT(13) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13]\, 
        F2H_INTERRUPT(12) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12]\, 
        F2H_INTERRUPT(11) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11]\, 
        F2H_INTERRUPT(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10]\, 
        F2H_INTERRUPT(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9]\, 
        F2H_INTERRUPT(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8]\, 
        F2H_INTERRUPT(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7]\, 
        F2H_INTERRUPT(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6]\, 
        F2H_INTERRUPT(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5]\, 
        F2H_INTERRUPT(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4]\, 
        F2H_INTERRUPT(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3]\, 
        F2H_INTERRUPT(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2]\, 
        F2H_INTERRUPT(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1]\, 
        F2H_INTERRUPT(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0]\, 
        F2HCALIB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2HCALIB_net\, 
        F_DMAREADY(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1]\, 
        F_DMAREADY(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0]\, 
        F_FM0_ADDR(31) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31]\, 
        F_FM0_ADDR(30) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30]\, 
        F_FM0_ADDR(29) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29]\, 
        F_FM0_ADDR(28) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28]\, 
        F_FM0_ADDR(27) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27]\, 
        F_FM0_ADDR(26) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26]\, 
        F_FM0_ADDR(25) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25]\, 
        F_FM0_ADDR(24) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24]\, 
        F_FM0_ADDR(23) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23]\, 
        F_FM0_ADDR(22) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22]\, 
        F_FM0_ADDR(21) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21]\, 
        F_FM0_ADDR(20) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20]\, 
        F_FM0_ADDR(19) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19]\, 
        F_FM0_ADDR(18) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18]\, 
        F_FM0_ADDR(17) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17]\, 
        F_FM0_ADDR(16) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16]\, 
        F_FM0_ADDR(15) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15]\, 
        F_FM0_ADDR(14) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14]\, 
        F_FM0_ADDR(13) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13]\, 
        F_FM0_ADDR(12) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12]\, 
        F_FM0_ADDR(11) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11]\, 
        F_FM0_ADDR(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10]\, 
        F_FM0_ADDR(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9]\, 
        F_FM0_ADDR(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8]\, 
        F_FM0_ADDR(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7]\, 
        F_FM0_ADDR(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6]\, 
        F_FM0_ADDR(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5]\, 
        F_FM0_ADDR(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4]\, 
        F_FM0_ADDR(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3]\, 
        F_FM0_ADDR(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2]\, 
        F_FM0_ADDR(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1]\, 
        F_FM0_ADDR(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0]\, 
        F_FM0_ENABLE => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net\, 
        F_FM0_MASTLOCK => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net\, 
        F_FM0_READY => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net\, 
        F_FM0_SEL => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net\, 
        F_FM0_SIZE(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1]\, 
        F_FM0_SIZE(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0]\, 
        F_FM0_TRANS1 => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net\, 
        F_FM0_WDATA(31) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31]\, 
        F_FM0_WDATA(30) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30]\, 
        F_FM0_WDATA(29) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29]\, 
        F_FM0_WDATA(28) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28]\, 
        F_FM0_WDATA(27) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27]\, 
        F_FM0_WDATA(26) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26]\, 
        F_FM0_WDATA(25) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25]\, 
        F_FM0_WDATA(24) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24]\, 
        F_FM0_WDATA(23) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23]\, 
        F_FM0_WDATA(22) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22]\, 
        F_FM0_WDATA(21) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21]\, 
        F_FM0_WDATA(20) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20]\, 
        F_FM0_WDATA(19) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19]\, 
        F_FM0_WDATA(18) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18]\, 
        F_FM0_WDATA(17) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17]\, 
        F_FM0_WDATA(16) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16]\, 
        F_FM0_WDATA(15) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15]\, 
        F_FM0_WDATA(14) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14]\, 
        F_FM0_WDATA(13) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13]\, 
        F_FM0_WDATA(12) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12]\, 
        F_FM0_WDATA(11) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11]\, 
        F_FM0_WDATA(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10]\, 
        F_FM0_WDATA(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9]\, 
        F_FM0_WDATA(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8]\, 
        F_FM0_WDATA(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7]\, 
        F_FM0_WDATA(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6]\, 
        F_FM0_WDATA(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5]\, 
        F_FM0_WDATA(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4]\, 
        F_FM0_WDATA(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3]\, 
        F_FM0_WDATA(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2]\, 
        F_FM0_WDATA(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1]\, 
        F_FM0_WDATA(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0]\, 
        F_FM0_WRITE => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net\, 
        F_HM0_RDATA(31) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31]\, 
        F_HM0_RDATA(30) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30]\, 
        F_HM0_RDATA(29) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29]\, 
        F_HM0_RDATA(28) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28]\, 
        F_HM0_RDATA(27) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27]\, 
        F_HM0_RDATA(26) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26]\, 
        F_HM0_RDATA(25) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25]\, 
        F_HM0_RDATA(24) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24]\, 
        F_HM0_RDATA(23) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23]\, 
        F_HM0_RDATA(22) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22]\, 
        F_HM0_RDATA(21) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21]\, 
        F_HM0_RDATA(20) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20]\, 
        F_HM0_RDATA(19) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19]\, 
        F_HM0_RDATA(18) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18]\, 
        F_HM0_RDATA(17) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17]\, 
        F_HM0_RDATA(16) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16]\, 
        F_HM0_RDATA(15) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15]\, 
        F_HM0_RDATA(14) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14]\, 
        F_HM0_RDATA(13) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13]\, 
        F_HM0_RDATA(12) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12]\, 
        F_HM0_RDATA(11) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11]\, 
        F_HM0_RDATA(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10]\, 
        F_HM0_RDATA(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9]\, 
        F_HM0_RDATA(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8]\, 
        F_HM0_RDATA(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7]\, 
        F_HM0_RDATA(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6]\, 
        F_HM0_RDATA(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5]\, 
        F_HM0_RDATA(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4]\, 
        F_HM0_RDATA(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3]\, 
        F_HM0_RDATA(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2]\, 
        F_HM0_RDATA(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1]\, 
        F_HM0_RDATA(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0]\, 
        F_HM0_READY => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net\, 
        F_HM0_RESP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net\, 
        FAB_AVALID => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net\, 
        FAB_HOSTDISCON => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net\, 
        FAB_IDDIG => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net\, 
        FAB_LINESTATE(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1]\, 
        FAB_LINESTATE(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0]\, 
        FAB_M3_RESET_N => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net\, 
        FAB_PLL_LOCK => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net\, 
        FAB_RXACTIVE => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net\, 
        FAB_RXERROR => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net\, 
        FAB_RXVALID => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net\, 
        FAB_RXVALIDH => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net\, 
        FAB_SESSEND => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net\, 
        FAB_TXREADY => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net\, 
        FAB_VBUSVALID => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net\, 
        FAB_VSTATUS(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7]\, 
        FAB_VSTATUS(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6]\, 
        FAB_VSTATUS(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5]\, 
        FAB_VSTATUS(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4]\, 
        FAB_VSTATUS(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3]\, 
        FAB_VSTATUS(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2]\, 
        FAB_VSTATUS(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1]\, 
        FAB_VSTATUS(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0]\, 
        FAB_XDATAIN(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7]\, 
        FAB_XDATAIN(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6]\, 
        FAB_XDATAIN(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5]\, 
        FAB_XDATAIN(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4]\, 
        FAB_XDATAIN(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3]\, 
        FAB_XDATAIN(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2]\, 
        FAB_XDATAIN(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1]\, 
        FAB_XDATAIN(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0]\, 
        GTX_CLKPF => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net\, 
        I2C0_BCLK => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net\, 
        I2C0_SCL_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net\, 
        I2C0_SDA_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net\, 
        I2C1_BCLK => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net\, 
        I2C1_SCL_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net\, 
        I2C1_SDA_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net\, 
        MDIF => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDIF_net\, 
        MGPIO0A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net\, 
        MGPIO10A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net\, 
        MGPIO11A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net\, 
        MGPIO11B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net\, 
        MGPIO12A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net\, 
        MGPIO13A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net\, 
        MGPIO14A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net\, 
        MGPIO15A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net\, 
        MGPIO16A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net\, 
        MGPIO17B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net\, 
        MGPIO18B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net\, 
        MGPIO19B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net\, 
        MGPIO1A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net\, 
        MGPIO20B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net\, 
        MGPIO21B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net\, 
        MGPIO22B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net\, 
        MGPIO24B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net\, 
        MGPIO25B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net\, 
        MGPIO26B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net\, 
        MGPIO27B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net\, 
        MGPIO28B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net\, 
        MGPIO29B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net\, 
        MGPIO2A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net\, 
        MGPIO30B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net\, 
        MGPIO31B_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net\, 
        MGPIO3A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net\, 
        MGPIO4A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net\, 
        MGPIO5A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net\, 
        MGPIO6A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net\, 
        MGPIO7A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net\, 
        MGPIO8A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net\, 
        MGPIO9A_F2H_GPIN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net\, 
        MMUART0_CTS_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net\, 
        MMUART0_DCD_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net\, 
        MMUART0_DSR_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net\, 
        MMUART0_DTR_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net\, 
        MMUART0_RI_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net\, 
        MMUART0_RTS_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net\, 
        MMUART0_RXD_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net\, 
        MMUART0_SCK_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net\, 
        MMUART0_TXD_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net\, 
        MMUART1_CTS_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net\, 
        MMUART1_DCD_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net\, 
        MMUART1_DSR_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net\, 
        MMUART1_RI_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net\, 
        MMUART1_RTS_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net\, 
        MMUART1_RXD_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net\, 
        MMUART1_SCK_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net\, 
        MMUART1_TXD_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net\, 
        PER2_FABRIC_PRDATA(31) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31]\, 
        PER2_FABRIC_PRDATA(30) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30]\, 
        PER2_FABRIC_PRDATA(29) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29]\, 
        PER2_FABRIC_PRDATA(28) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28]\, 
        PER2_FABRIC_PRDATA(27) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27]\, 
        PER2_FABRIC_PRDATA(26) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26]\, 
        PER2_FABRIC_PRDATA(25) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25]\, 
        PER2_FABRIC_PRDATA(24) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24]\, 
        PER2_FABRIC_PRDATA(23) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23]\, 
        PER2_FABRIC_PRDATA(22) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22]\, 
        PER2_FABRIC_PRDATA(21) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21]\, 
        PER2_FABRIC_PRDATA(20) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20]\, 
        PER2_FABRIC_PRDATA(19) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19]\, 
        PER2_FABRIC_PRDATA(18) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18]\, 
        PER2_FABRIC_PRDATA(17) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17]\, 
        PER2_FABRIC_PRDATA(16) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16]\, 
        PER2_FABRIC_PRDATA(15) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15]\, 
        PER2_FABRIC_PRDATA(14) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14]\, 
        PER2_FABRIC_PRDATA(13) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13]\, 
        PER2_FABRIC_PRDATA(12) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12]\, 
        PER2_FABRIC_PRDATA(11) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11]\, 
        PER2_FABRIC_PRDATA(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10]\, 
        PER2_FABRIC_PRDATA(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9]\, 
        PER2_FABRIC_PRDATA(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8]\, 
        PER2_FABRIC_PRDATA(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7]\, 
        PER2_FABRIC_PRDATA(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6]\, 
        PER2_FABRIC_PRDATA(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5]\, 
        PER2_FABRIC_PRDATA(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4]\, 
        PER2_FABRIC_PRDATA(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3]\, 
        PER2_FABRIC_PRDATA(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2]\, 
        PER2_FABRIC_PRDATA(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1]\, 
        PER2_FABRIC_PRDATA(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0]\, 
        PER2_FABRIC_PREADY => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net\, 
        PER2_FABRIC_PSLVERR => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net\, 
        RCGF(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[9]\, RCGF(8)
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[8]\, 
        RCGF(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[7]\, RCGF(6)
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[6]\, 
        RCGF(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[5]\, RCGF(4)
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[4]\, 
        RCGF(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[3]\, RCGF(2)
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[2]\, 
        RCGF(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[1]\, RCGF(0)
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[0]\, 
        RX_CLKPF => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net\, RX_DVF
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_DVF_net\, 
        RX_ERRF => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_ERRF_net\, RX_EV
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_EV_net\, 
        RXDF(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[7]\, RXDF(6)
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[6]\, 
        RXDF(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[5]\, RXDF(4)
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[4]\, 
        RXDF(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[3]\, RXDF(2)
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[2]\, 
        RXDF(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[1]\, RXDF(0)
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[0]\, 
        SLEEPHOLDREQ => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net\, 
        SMBALERT_NI0 => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net\, 
        SMBALERT_NI1 => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net\, 
        SMBSUS_NI0 => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net\, 
        SMBSUS_NI1 => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net\, 
        SPI0_CLK_IN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net\, 
        SPI0_SDI_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net\, 
        SPI0_SDO_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net\, 
        SPI0_SS0_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net\, 
        SPI0_SS1_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net\, 
        SPI0_SS2_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net\, 
        SPI0_SS3_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net\, 
        SPI1_CLK_IN => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net\, 
        SPI1_SDI_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net\, 
        SPI1_SDO_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net\, 
        SPI1_SS0_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net\, 
        SPI1_SS1_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net\, 
        SPI1_SS2_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net\, 
        SPI1_SS3_F2H_SCP => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net\, 
        TX_CLKPF => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net\, 
        USER_MSS_GPIO_RESET_N => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net\, 
        USER_MSS_RESET_N => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net\, 
        XCLK_FAB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net\, 
        CLK_BASE => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CLK_BASE_net\, 
        CLK_MDDR_APB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net\, 
        F_ARADDR_HADDR1(31) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31]\, 
        F_ARADDR_HADDR1(30) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30]\, 
        F_ARADDR_HADDR1(29) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29]\, 
        F_ARADDR_HADDR1(28) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28]\, 
        F_ARADDR_HADDR1(27) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27]\, 
        F_ARADDR_HADDR1(26) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26]\, 
        F_ARADDR_HADDR1(25) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25]\, 
        F_ARADDR_HADDR1(24) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24]\, 
        F_ARADDR_HADDR1(23) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23]\, 
        F_ARADDR_HADDR1(22) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22]\, 
        F_ARADDR_HADDR1(21) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21]\, 
        F_ARADDR_HADDR1(20) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20]\, 
        F_ARADDR_HADDR1(19) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19]\, 
        F_ARADDR_HADDR1(18) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18]\, 
        F_ARADDR_HADDR1(17) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17]\, 
        F_ARADDR_HADDR1(16) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16]\, 
        F_ARADDR_HADDR1(15) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15]\, 
        F_ARADDR_HADDR1(14) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14]\, 
        F_ARADDR_HADDR1(13) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13]\, 
        F_ARADDR_HADDR1(12) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12]\, 
        F_ARADDR_HADDR1(11) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11]\, 
        F_ARADDR_HADDR1(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10]\, 
        F_ARADDR_HADDR1(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9]\, 
        F_ARADDR_HADDR1(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8]\, 
        F_ARADDR_HADDR1(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7]\, 
        F_ARADDR_HADDR1(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6]\, 
        F_ARADDR_HADDR1(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5]\, 
        F_ARADDR_HADDR1(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4]\, 
        F_ARADDR_HADDR1(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3]\, 
        F_ARADDR_HADDR1(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2]\, 
        F_ARADDR_HADDR1(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1]\, 
        F_ARADDR_HADDR1(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0]\, 
        F_ARBURST_HTRANS1(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1]\, 
        F_ARBURST_HTRANS1(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0]\, 
        F_ARID_HSEL1(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3]\, 
        F_ARID_HSEL1(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2]\, 
        F_ARID_HSEL1(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1]\, 
        F_ARID_HSEL1(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0]\, 
        F_ARLEN_HBURST1(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3]\, 
        F_ARLEN_HBURST1(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2]\, 
        F_ARLEN_HBURST1(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1]\, 
        F_ARLEN_HBURST1(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0]\, 
        F_ARLOCK_HMASTLOCK1(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1]\, 
        F_ARLOCK_HMASTLOCK1(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0]\, 
        F_ARSIZE_HSIZE1(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1]\, 
        F_ARSIZE_HSIZE1(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0]\, 
        F_ARVALID_HWRITE1 => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net\, 
        F_AWADDR_HADDR0(31) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31]\, 
        F_AWADDR_HADDR0(30) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30]\, 
        F_AWADDR_HADDR0(29) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29]\, 
        F_AWADDR_HADDR0(28) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28]\, 
        F_AWADDR_HADDR0(27) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27]\, 
        F_AWADDR_HADDR0(26) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26]\, 
        F_AWADDR_HADDR0(25) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25]\, 
        F_AWADDR_HADDR0(24) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24]\, 
        F_AWADDR_HADDR0(23) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23]\, 
        F_AWADDR_HADDR0(22) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22]\, 
        F_AWADDR_HADDR0(21) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21]\, 
        F_AWADDR_HADDR0(20) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20]\, 
        F_AWADDR_HADDR0(19) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19]\, 
        F_AWADDR_HADDR0(18) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18]\, 
        F_AWADDR_HADDR0(17) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17]\, 
        F_AWADDR_HADDR0(16) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16]\, 
        F_AWADDR_HADDR0(15) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15]\, 
        F_AWADDR_HADDR0(14) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14]\, 
        F_AWADDR_HADDR0(13) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13]\, 
        F_AWADDR_HADDR0(12) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12]\, 
        F_AWADDR_HADDR0(11) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11]\, 
        F_AWADDR_HADDR0(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10]\, 
        F_AWADDR_HADDR0(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9]\, 
        F_AWADDR_HADDR0(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8]\, 
        F_AWADDR_HADDR0(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7]\, 
        F_AWADDR_HADDR0(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6]\, 
        F_AWADDR_HADDR0(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5]\, 
        F_AWADDR_HADDR0(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4]\, 
        F_AWADDR_HADDR0(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3]\, 
        F_AWADDR_HADDR0(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2]\, 
        F_AWADDR_HADDR0(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1]\, 
        F_AWADDR_HADDR0(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0]\, 
        F_AWBURST_HTRANS0(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1]\, 
        F_AWBURST_HTRANS0(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0]\, 
        F_AWID_HSEL0(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3]\, 
        F_AWID_HSEL0(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2]\, 
        F_AWID_HSEL0(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1]\, 
        F_AWID_HSEL0(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0]\, 
        F_AWLEN_HBURST0(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3]\, 
        F_AWLEN_HBURST0(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2]\, 
        F_AWLEN_HBURST0(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1]\, 
        F_AWLEN_HBURST0(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0]\, 
        F_AWLOCK_HMASTLOCK0(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1]\, 
        F_AWLOCK_HMASTLOCK0(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0]\, 
        F_AWSIZE_HSIZE0(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1]\, 
        F_AWSIZE_HSIZE0(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0]\, 
        F_AWVALID_HWRITE0 => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net\, 
        F_BREADY => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_BREADY_net\, 
        F_RMW_AXI => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net\, 
        F_RREADY => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_RREADY_net\, 
        F_WDATA_HWDATA01(63) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63]\, 
        F_WDATA_HWDATA01(62) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62]\, 
        F_WDATA_HWDATA01(61) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61]\, 
        F_WDATA_HWDATA01(60) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60]\, 
        F_WDATA_HWDATA01(59) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59]\, 
        F_WDATA_HWDATA01(58) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58]\, 
        F_WDATA_HWDATA01(57) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57]\, 
        F_WDATA_HWDATA01(56) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56]\, 
        F_WDATA_HWDATA01(55) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55]\, 
        F_WDATA_HWDATA01(54) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54]\, 
        F_WDATA_HWDATA01(53) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53]\, 
        F_WDATA_HWDATA01(52) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52]\, 
        F_WDATA_HWDATA01(51) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51]\, 
        F_WDATA_HWDATA01(50) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50]\, 
        F_WDATA_HWDATA01(49) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49]\, 
        F_WDATA_HWDATA01(48) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48]\, 
        F_WDATA_HWDATA01(47) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47]\, 
        F_WDATA_HWDATA01(46) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46]\, 
        F_WDATA_HWDATA01(45) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45]\, 
        F_WDATA_HWDATA01(44) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44]\, 
        F_WDATA_HWDATA01(43) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43]\, 
        F_WDATA_HWDATA01(42) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42]\, 
        F_WDATA_HWDATA01(41) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41]\, 
        F_WDATA_HWDATA01(40) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40]\, 
        F_WDATA_HWDATA01(39) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39]\, 
        F_WDATA_HWDATA01(38) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38]\, 
        F_WDATA_HWDATA01(37) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37]\, 
        F_WDATA_HWDATA01(36) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36]\, 
        F_WDATA_HWDATA01(35) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35]\, 
        F_WDATA_HWDATA01(34) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34]\, 
        F_WDATA_HWDATA01(33) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33]\, 
        F_WDATA_HWDATA01(32) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32]\, 
        F_WDATA_HWDATA01(31) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31]\, 
        F_WDATA_HWDATA01(30) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30]\, 
        F_WDATA_HWDATA01(29) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29]\, 
        F_WDATA_HWDATA01(28) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28]\, 
        F_WDATA_HWDATA01(27) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27]\, 
        F_WDATA_HWDATA01(26) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26]\, 
        F_WDATA_HWDATA01(25) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25]\, 
        F_WDATA_HWDATA01(24) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24]\, 
        F_WDATA_HWDATA01(23) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23]\, 
        F_WDATA_HWDATA01(22) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22]\, 
        F_WDATA_HWDATA01(21) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21]\, 
        F_WDATA_HWDATA01(20) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20]\, 
        F_WDATA_HWDATA01(19) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19]\, 
        F_WDATA_HWDATA01(18) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18]\, 
        F_WDATA_HWDATA01(17) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17]\, 
        F_WDATA_HWDATA01(16) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16]\, 
        F_WDATA_HWDATA01(15) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15]\, 
        F_WDATA_HWDATA01(14) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14]\, 
        F_WDATA_HWDATA01(13) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13]\, 
        F_WDATA_HWDATA01(12) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12]\, 
        F_WDATA_HWDATA01(11) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11]\, 
        F_WDATA_HWDATA01(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10]\, 
        F_WDATA_HWDATA01(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9]\, 
        F_WDATA_HWDATA01(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8]\, 
        F_WDATA_HWDATA01(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7]\, 
        F_WDATA_HWDATA01(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6]\, 
        F_WDATA_HWDATA01(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5]\, 
        F_WDATA_HWDATA01(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4]\, 
        F_WDATA_HWDATA01(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3]\, 
        F_WDATA_HWDATA01(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2]\, 
        F_WDATA_HWDATA01(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1]\, 
        F_WDATA_HWDATA01(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0]\, 
        F_WID_HREADY01(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3]\, 
        F_WID_HREADY01(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2]\, 
        F_WID_HREADY01(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1]\, 
        F_WID_HREADY01(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0]\, 
        F_WLAST => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WLAST_net\, 
        F_WSTRB(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7]\, 
        F_WSTRB(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6]\, 
        F_WSTRB(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5]\, 
        F_WSTRB(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4]\, 
        F_WSTRB(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3]\, 
        F_WSTRB(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2]\, 
        F_WSTRB(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1]\, 
        F_WSTRB(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0]\, 
        F_WVALID => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WVALID_net\, 
        FPGA_MDDR_ARESET_N => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net\, 
        MDDR_FABRIC_PADDR(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10]\, 
        MDDR_FABRIC_PADDR(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9]\, 
        MDDR_FABRIC_PADDR(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8]\, 
        MDDR_FABRIC_PADDR(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7]\, 
        MDDR_FABRIC_PADDR(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6]\, 
        MDDR_FABRIC_PADDR(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5]\, 
        MDDR_FABRIC_PADDR(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4]\, 
        MDDR_FABRIC_PADDR(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3]\, 
        MDDR_FABRIC_PADDR(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2]\, 
        MDDR_FABRIC_PENABLE => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net\, 
        MDDR_FABRIC_PSEL => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net\, 
        MDDR_FABRIC_PWDATA(15) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15]\, 
        MDDR_FABRIC_PWDATA(14) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14]\, 
        MDDR_FABRIC_PWDATA(13) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13]\, 
        MDDR_FABRIC_PWDATA(12) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12]\, 
        MDDR_FABRIC_PWDATA(11) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11]\, 
        MDDR_FABRIC_PWDATA(10) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10]\, 
        MDDR_FABRIC_PWDATA(9) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9]\, 
        MDDR_FABRIC_PWDATA(8) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8]\, 
        MDDR_FABRIC_PWDATA(7) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7]\, 
        MDDR_FABRIC_PWDATA(6) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6]\, 
        MDDR_FABRIC_PWDATA(5) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5]\, 
        MDDR_FABRIC_PWDATA(4) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4]\, 
        MDDR_FABRIC_PWDATA(3) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3]\, 
        MDDR_FABRIC_PWDATA(2) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2]\, 
        MDDR_FABRIC_PWDATA(1) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1]\, 
        MDDR_FABRIC_PWDATA(0) => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0]\, 
        MDDR_FABRIC_PWRITE => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net\, 
        PRESET_N => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PRESET_N_net\, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => ADLIB_GND0, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => ADLIB_GND0, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => ADLIB_GND0, DM_IN(2)
         => ADLIB_GND0, DM_IN(1) => ADLIB_GND0, DM_IN(0) => 
        ADLIB_GND0, DRAM_DQ_IN(17) => ADLIB_GND0, DRAM_DQ_IN(16)
         => ADLIB_GND0, DRAM_DQ_IN(15) => ADLIB_GND0, 
        DRAM_DQ_IN(14) => ADLIB_GND0, DRAM_DQ_IN(13) => 
        ADLIB_GND0, DRAM_DQ_IN(12) => ADLIB_GND0, DRAM_DQ_IN(11)
         => ADLIB_GND0, DRAM_DQ_IN(10) => ADLIB_GND0, 
        DRAM_DQ_IN(9) => ADLIB_GND0, DRAM_DQ_IN(8) => ADLIB_GND0, 
        DRAM_DQ_IN(7) => ADLIB_GND0, DRAM_DQ_IN(6) => ADLIB_GND0, 
        DRAM_DQ_IN(5) => ADLIB_GND0, DRAM_DQ_IN(4) => ADLIB_GND0, 
        DRAM_DQ_IN(3) => ADLIB_GND0, DRAM_DQ_IN(2) => ADLIB_GND0, 
        DRAM_DQ_IN(1) => ADLIB_GND0, DRAM_DQ_IN(0) => ADLIB_GND0, 
        DRAM_DQS_IN(2) => ADLIB_GND0, DRAM_DQS_IN(1) => 
        ADLIB_GND0, DRAM_DQS_IN(0) => ADLIB_GND0, 
        DRAM_FIFO_WE_IN(1) => ADLIB_GND0, DRAM_FIFO_WE_IN(0) => 
        ADLIB_GND0, I2C0_SCL_USBC_DATA1_MGPIO31B_IN => ADLIB_GND0, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => ADLIB_GND0, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => ADLIB_GND0, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => ADLIB_GND0, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => ADLIB_GND0, 
        MMUART0_DCD_MGPIO22B_IN => ADLIB_GND0, 
        MMUART0_DSR_MGPIO20B_IN => ADLIB_GND0, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => ADLIB_GND0, 
        MMUART0_RI_MGPIO21B_IN => ADLIB_GND0, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => ADLIB_GND0, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => ADLIB_GND0, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => ADLIB_GND0, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => ADLIB_GND0, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => ADLIB_GND0, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => ADLIB_GND0, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => ADLIB_GND0, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => ADLIB_GND0, 
        RGMII_MDC_RMII_MDC_IN => ADLIB_GND0, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => ADLIB_GND0, 
        RGMII_RX_CLK_IN => ADLIB_GND0, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => ADLIB_GND0, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => ADLIB_GND0, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => ADLIB_GND0, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => ADLIB_GND0, 
        RGMII_RXD3_USBB_DATA4_IN => ADLIB_GND0, RGMII_TX_CLK_IN
         => ADLIB_GND0, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        ADLIB_GND0, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => 
        ADLIB_GND0, RGMII_TXD1_RMII_TXD1_USBB_STP_IN => 
        ADLIB_GND0, RGMII_TXD2_USBB_DATA5_IN => ADLIB_GND0, 
        RGMII_TXD3_USBB_DATA6_IN => ADLIB_GND0, 
        SPI0_SCK_USBA_XCLK_IN => ADLIB_GND0, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => ADLIB_GND0, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => ADLIB_GND0, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => ADLIB_GND0, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => ADLIB_GND0, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => ADLIB_GND0, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => ADLIB_GND0, 
        SPI1_SCK_IN => ADLIB_GND0, SPI1_SDI_MGPIO11A_IN => 
        ADLIB_GND0, SPI1_SDO_MGPIO12A_IN => ADLIB_GND0, 
        SPI1_SS0_MGPIO13A_IN => ADLIB_GND0, SPI1_SS1_MGPIO14A_IN
         => ADLIB_GND0, SPI1_SS2_MGPIO15A_IN => ADLIB_GND0, 
        SPI1_SS3_MGPIO16A_IN => ADLIB_GND0, SPI1_SS4_MGPIO17A_IN
         => ADLIB_GND0, SPI1_SS5_MGPIO18A_IN => ADLIB_GND0, 
        SPI1_SS6_MGPIO23A_IN => ADLIB_GND0, SPI1_SS7_MGPIO24A_IN
         => ADLIB_GND0, USBC_XCLK_IN => ADLIB_GND0, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => nc239, DRAM_ADDR(14) => nc353, DRAM_ADDR(13) => nc348, 
        DRAM_ADDR(12) => nc142, DRAM_ADDR(11) => nc320, 
        DRAM_ADDR(10) => nc344, DRAM_ADDR(9) => nc315, 
        DRAM_ADDR(8) => nc382, DRAM_ADDR(7) => nc247, 
        DRAM_ADDR(6) => nc94, DRAM_ADDR(5) => nc197, DRAM_ADDR(4)
         => nc328, DRAM_ADDR(3) => nc122, DRAM_ADDR(2) => nc266, 
        DRAM_ADDR(1) => nc35, DRAM_ADDR(0) => nc324, DRAM_BA(2)
         => nc4, DRAM_BA(1) => nc227, DRAM_BA(0) => nc92, 
        DRAM_CASN => OPEN, DRAM_CKE => OPEN, DRAM_CLK => OPEN, 
        DRAM_CSN => OPEN, DRAM_DM_RDQS_OUT(2) => nc101, 
        DRAM_DM_RDQS_OUT(1) => nc413, DRAM_DM_RDQS_OUT(0) => 
        nc346, DRAM_DQ_OUT(17) => nc330, DRAM_DQ_OUT(16) => nc397, 
        DRAM_DQ_OUT(15) => nc184, DRAM_DQ_OUT(14) => nc200, 
        DRAM_DQ_OUT(13) => nc190, DRAM_DQ_OUT(12) => nc166, 
        DRAM_DQ_OUT(11) => nc372, DRAM_DQ_OUT(10) => nc407, 
        DRAM_DQ_OUT(9) => nc355, DRAM_DQ_OUT(8) => nc338, 
        DRAM_DQ_OUT(7) => nc326, DRAM_DQ_OUT(6) => nc132, 
        DRAM_DQ_OUT(5) => nc383, DRAM_DQ_OUT(4) => nc334, 
        DRAM_DQ_OUT(3) => nc21, DRAM_DQ_OUT(2) => nc237, 
        DRAM_DQ_OUT(1) => nc93, DRAM_DQ_OUT(0) => nc262, 
        DRAM_DQS_OUT(2) => nc69, DRAM_DQS_OUT(1) => nc206, 
        DRAM_DQS_OUT(0) => nc174, DRAM_FIFO_WE_OUT(1) => nc38, 
        DRAM_FIFO_WE_OUT(0) => nc113, DRAM_ODT => OPEN, DRAM_RASN
         => OPEN, DRAM_RSTN => OPEN, DRAM_WEN => OPEN, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OUT => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT => OPEN, 
        MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => OPEN, SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, SPI1_SCK_OUT
         => OPEN, SPI1_SDI_MGPIO11A_OUT => OPEN, 
        SPI1_SDO_MGPIO12A_OUT => OPEN, SPI1_SS0_MGPIO13A_OUT => 
        OPEN, SPI1_SS1_MGPIO14A_OUT => OPEN, 
        SPI1_SS2_MGPIO15A_OUT => OPEN, SPI1_SS3_MGPIO16A_OUT => 
        OPEN, SPI1_SS4_MGPIO17A_OUT => OPEN, 
        SPI1_SS5_MGPIO18A_OUT => OPEN, SPI1_SS6_MGPIO23A_OUT => 
        OPEN, SPI1_SS7_MGPIO24A_OUT => OPEN, USBC_XCLK_OUT => 
        OPEN, CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => OPEN, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => 
        nc336, DM_OE(1) => nc218, DM_OE(0) => nc401, 
        DRAM_DQ_OE(17) => nc342, DRAM_DQ_OE(16) => nc373, 
        DRAM_DQ_OE(15) => nc106, DRAM_DQ_OE(14) => nc261, 
        DRAM_DQ_OE(13) => nc25, DRAM_DQ_OE(12) => nc1, 
        DRAM_DQ_OE(11) => nc385, DRAM_DQ_OE(10) => nc426, 
        DRAM_DQ_OE(9) => nc322, DRAM_DQ_OE(8) => nc299, 
        DRAM_DQ_OE(7) => nc37, DRAM_DQ_OE(6) => nc410, 
        DRAM_DQ_OE(5) => nc202, DRAM_DQ_OE(4) => nc144, 
        DRAM_DQ_OE(3) => nc153, DRAM_DQ_OE(2) => nc46, 
        DRAM_DQ_OE(1) => nc258, DRAM_DQ_OE(0) => nc343, 
        DRAM_DQS_OE(2) => nc71, DRAM_DQS_OE(1) => nc124, 
        DRAM_DQS_OE(0) => nc436, I2C0_SCL_USBC_DATA1_MGPIO31B_OE
         => OPEN, I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => OPEN, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => OPEN, SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => OPEN, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => OPEN, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => OPEN, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, SPI1_SCK_OE => 
        OPEN, SPI1_SDI_MGPIO11A_OE => OPEN, SPI1_SDO_MGPIO12A_OE
         => OPEN, SPI1_SS0_MGPIO13A_OE => OPEN, 
        SPI1_SS1_MGPIO14A_OE => OPEN, SPI1_SS2_MGPIO15A_OE => 
        OPEN, SPI1_SS3_MGPIO16A_OE => OPEN, SPI1_SS4_MGPIO17A_OE
         => OPEN, SPI1_SS5_MGPIO18A_OE => OPEN, 
        SPI1_SS6_MGPIO23A_OE => OPEN, SPI1_SS7_MGPIO24A_OE => 
        OPEN, USBC_XCLK_OE => OPEN);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[9]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[9]\, B => 
        \sb_sb_0_Memory_PRDATA[9]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9]\);
    
    \MemorySynchronizer_0/SynchStatusReg_152_e2_0_a2_0_a2\ : CFG3
      generic map(INIT => x"02")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[2]\, 
        B => \MemorySynchronizer_0/MemorySyncState_Z[3]\, C => 
        \MemorySynchronizer_0/un1_enabletimestampgen2_2_sn\, Y
         => \MemorySynchronizer_0/SynchStatusReg_152_e2\);
    
    \STAMP_0/spi/rx_data[10]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[10]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_39_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_59\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_39_set_Z\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[6]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[6]\);
    
    \MemorySynchronizer_0/un1_nreset_57_0_a3_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[9]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_57_i\);
    
    \STAMP_0/spi/un7_count_NE_20_RNIK2531\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \STAMP_0/spi/un7_count_NE_20_Z\, B => 
        \STAMP_0/spi/un7_count_NE_21_Z\, C => 
        \STAMP_0/spi/un7_count_NE_28_Z\, D => 
        \STAMP_0/spi/un7_count_NE_27_Z\, Y => 
        \STAMP_0/spi/un7_count_NE_i\);
    
    \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_3_i_0_a2_0\ : 
        CFG3
      generic map(INIT => x"08")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_2561\, C => 
        \sb_sb_0_STAMP_PADDR[4]\, Y => 
        \MemorySynchronizer_0/N_2517\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_38\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[2]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[2]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1089\, Y => 
        \MemorySynchronizer_0/N_1120\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[22]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[22]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[10]\, Y
         => \MemorySynchronizer_0/N_1069\);
    
    \STAMP_0/dummy[13]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_60\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[13]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[18]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[18]\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/N_2323\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[18]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[18]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_211\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_43_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_61\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_43_set_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[1]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[1]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[1]\, C => 
        \MemorySynchronizer_0/N_2596\, D => 
        \MemorySynchronizer_0/N_2595\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[1]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[0]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[0]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[0]\, D => 
        \MemorySynchronizer_0/un5_resettimercounter_m[32]\, Y => 
        \MemorySynchronizer_0/resettimercounter_9[0]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_174\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net\, 
        IPC => OPEN);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_12\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/NGMUX0_ARST_N_net\, IPB
         => OPEN, IPC => \sb_sb_0/CCC_0/CCC_INST/PADDR_net[2]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[0]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[0]\);
    
    \STAMP_0/spi/rx_data[12]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[12]\);
    
    \STAMP_0/un1_spi_rx_data_2[18]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_601\, B => \STAMP_0/N_635\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_668\);
    
    \MemorySynchronizer_0/un1_in_enable_2_0_0_a2_0\ : CFG4
      generic map(INIT => x"0700")

      port map(A => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_28_Z\, 
        B => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_29_Z\, 
        C => STAMP_0_new_avail, D => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[15]\, Y
         => \MemorySynchronizer_0/N_2604\);
    
    \STAMP_0/spi_tx_data_RNO[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[7]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_291_i\);
    
    \MemorySynchronizer_0/un1_nreset_8_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_34_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_8_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_8_rs_Z\);
    
    \STAMP_0/dummy[5]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_62\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[5]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[15]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[15]\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2564\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1453\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_39_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[21]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_39\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_0[4]\ : 
        CFG4
      generic map(INIT => x"3320")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_2_0_Z[4]\, 
        B => STAMP_0_new_avail, C => 
        \MemorySynchronizer_0/N_2310\, D => 
        \MemorySynchronizer_0/N_1512\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_0_Z[4]\);
    
    \stamp0_spi_dms2_cs_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => stamp0_spi_dms2_cs_c, E => ADLIB_VCC1, DOUT
         => \stamp0_spi_dms2_cs_obuf/U0/DOUT1\, EOUT => 
        \stamp0_spi_dms2_cs_obuf/U0/EOUT1\);
    
    \STAMP_0/measurement_dms2[2]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[34]\);
    
    \MemorySynchronizer_0/un1_nreset_22_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_40\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_22_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_22_rs_Z\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[29]\ : SLE
      port map(D => \STAMP_0_data_frame[29]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[29]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[11]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[11]\);
    
    \stamp0_ready_temp_ibuf/U0/U_IOPAD\ : sdf_IOPAD_IN
      port map(PAD => stamp0_ready_temp, Y => 
        \stamp0_ready_temp_ibuf/U0/YIN1\);
    
    \STAMP_0/delay_counter_cry[10]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[10]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[9]\, S
         => \STAMP_0/delay_counter_s[10]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[10]\, CC => NET_CC_CONFIG425, 
        P => NET_CC_CONFIG423, UB => NET_CC_CONFIG424);
    
    AFLSDF_INV_24 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_42_Z\, Y => 
        \AFLSDF_INV_24\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[0]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[0]\, 
        B => \sb_sb_0_STAMP_PWDATA[0]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[0]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1[31]\ : 
        CFG4
      generic map(INIT => x"7FFF")

      port map(A => \MemorySynchronizer_0/N_2567\, B => 
        \MemorySynchronizer_0/N_2561\, C => 
        \MemorySynchronizer_0/APBState_Z[0]\, D => 
        \sb_sb_0_STAMP_PADDR[6]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_4\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX0_HOLD_N_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[2]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[1]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[1]\);
    
    AFLSDF_INV_84 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_34_Z\, Y => 
        \AFLSDF_INV_84\);
    
    \MemorySynchronizer_0/resynctimercounter[2]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1120\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[2]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_93\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RX_DVF_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_25\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[25]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_24_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[25]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_25_Z\, 
        CC => NET_CC_CONFIG179, P => NET_CC_CONFIG177, UB => 
        NET_CC_CONFIG178);
    
    \STAMP_0/spi/count_lm_0[27]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[27]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[27]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[23]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[23]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1068\, Y => 
        \MemorySynchronizer_0/N_1099\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[22]\ : SLE
      port map(D => \STAMP_0_data_frame[54]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[22]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_203\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19]\, 
        IPC => OPEN);
    
    AFLSDF_INV_50 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_38\, Y => 
        \AFLSDF_INV_50\);
    
    \MemorySynchronizer_0/SynchStatusReg2_RNO[21]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \MemorySynchronizer_0/temp_1_cry_0_Y\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[21]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[21]\);
    
    \MemorySynchronizer_0/PRDATA[6]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[6]\);
    
    \STAMP_0/spi_tx_data[2]\ : SLE
      port map(D => \STAMP_0/N_296_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[2]\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_63\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[21]\, B => 
        \MemorySynchronizer_0/un104_in_enable_20\, C => 
        \MemorySynchronizer_0/un104_in_enable_21\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[20]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[9]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[10]\, CC
         => NET_CC_CONFIG568, P => NET_CC_CONFIG566, UB => 
        NET_CC_CONFIG567);
    
    \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0\ : CFG4
      generic map(INIT => x"FDCC")

      port map(A => \MemorySynchronizer_0/N_140_2\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_0_Z\, 
        C => \MemorySynchronizer_0/SynchStatusReg_N_3_mux\, D => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_1_Z\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[12]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[12]\);
    
    \STAMP_0/dummy[2]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_63\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[2]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[13]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[13]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_43_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_64\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_43_set_Z\);
    
    \STAMP_0/spi/clk_toggles_s_390\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/spi/clk_toggles_Z[0]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => ADLIB_VCC1, S => OPEN, Y => OPEN, FCO
         => \STAMP_0/spi/clk_toggles_s_390_FCO\, CC => 
        NET_CC_CONFIG607, P => NET_CC_CONFIG605, UB => 
        NET_CC_CONFIG606);
    
    \MemorySynchronizer_0/ConfigReg[5]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[5]\);
    
    \STAMP_0/un1_spi_rx_data_0[14]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[14]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[14]\, Y
         => \STAMP_0/N_597\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[22]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[22]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[22]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[22]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[22]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[22]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_5\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[5]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_4_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_5_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_5_Z\, CC
         => NET_CC_CONFIG740, P => NET_CC_CONFIG738, UB => 
        NET_CC_CONFIG739);
    
    \STAMP_0/un1_PREADY_0_sqmuxa_3_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \STAMP_0/component_state_Z[4]\, B => 
        \STAMP_0/component_state_Z[5]\, C => \STAMP_0/N_162_i\, D
         => \STAMP_0/PREADY_0_sqmuxa_2\, Y => 
        \STAMP_0/un1_PREADY_0_sqmuxa_3_0_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg2[8]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[8]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[8]\);
    
    \STAMP_0/delay_counter[14]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[14]\);
    
    \STAMP_0/component_state_ns_0_0_0[2]\ : CFG4
      generic map(INIT => x"AEAA")

      port map(A => \STAMP_0/apb_spi_finished_0_sqmuxa\, B => 
        \STAMP_0/component_state_ns_0_0_a3_1_Z[2]\, C => 
        \STAMP_0/un27_paddr_i_0\, D => \STAMP_0/un13_paddr_i_0\, 
        Y => \STAMP_0/component_state_ns_0_0_0_Z[2]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_0_iv_0_0[31]\ : 
        CFG4
      generic map(INIT => x"CCEC")

      port map(A => \MemorySynchronizer_0/N_140_i\, B => 
        \MemorySynchronizer_0/N_2471\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_s_31_S\, 
        D => \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, 
        Y => \MemorySynchronizer_0/waitingtimercounter_10[31]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_1\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_2\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_0_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[2]\, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_1_Z\, 
        CC => NET_CC_CONFIG1026, P => NET_CC_CONFIG1024, UB => 
        NET_CC_CONFIG1025);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_7\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_8\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_6_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[8]\, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_7_Z\, 
        CC => NET_CC_CONFIG1044, P => NET_CC_CONFIG1042, UB => 
        NET_CC_CONFIG1043);
    
    \STAMP_0/un1_drdy_flank_detected_dms1_0_sqmuxa_1\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/un1_new_avail_0_sqmuxa_1\, B => 
        \STAMP_0/drdy_flank_detected_dms1_0_sqmuxa_1\, Y => 
        \STAMP_0/un1_drdy_flank_detected_dms1_0_sqmuxa_1_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_120\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/spi/count[12]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[12]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_102\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[2]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[9]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_27\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[27]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_26_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[27]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_27_Z\, 
        CC => NET_CC_CONFIG185, P => NET_CC_CONFIG183, UB => 
        NET_CC_CONFIG184);
    
    \STAMP_0/delay_counter_lm_0[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_216_i\, B => 
        \STAMP_0/component_state_RNIFR114_Z[0]\, C => 
        \STAMP_0/delay_counter_s[4]\, Y => 
        \STAMP_0/delay_counter_lm[4]\);
    
    \STAMP_0/spi/rx_data[7]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[7]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[25]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[25]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[24]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[25]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[25]\, CC
         => NET_CC_CONFIG81, P => NET_CC_CONFIG79, UB => 
        NET_CC_CONFIG80);
    
    \MemorySynchronizer_0/un1_nreset_4_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[4]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_4_i\);
    
    \MemorySynchronizer_0/un1_MemorySyncState_11\ : CFG4
      generic map(INIT => x"CEEE")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => \MemorySynchronizer_0/MemorySyncState_Z[5]\, C => 
        \MemorySynchronizer_0/un94_in_enable_29_Z\, D => 
        \MemorySynchronizer_0/un94_in_enable_28_Z\, Y => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\);
    
    \MemorySynchronizer_0/N_1980_i_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_65\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_1980_i_set_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[1]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_1\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[1]\, 
        C => \MemorySynchronizer_0/N_1561\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[1]\);
    
    \stamp0_ready_dms1_ibuf/U0/U_IOINFF\ : IOINFF_BYPASS
      port map(A => \stamp0_ready_dms1_ibuf/U0/YIN1\, Y => 
        \stamp0_ready_dms1_ibuf/U0/YIN\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[13]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[13]\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_13_S\, 
        C => \MemorySynchronizer_0/resettimercounter_m[13]\, D
         => \MemorySynchronizer_0/resettimercounter_0_sqmuxa_1\, 
        Y => \MemorySynchronizer_0/resettimercounter_9[13]\);
    
    \MemorySynchronizer_0/un1_nreset_29\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[25]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_29_i\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[20]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[20]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[20]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[20]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_16\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[16]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[16]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_15_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_16_Z\, CC => 
        NET_CC_CONFIG871, P => NET_CC_CONFIG869, UB => 
        NET_CC_CONFIG870);
    
    \MemorySynchronizer_0/SynchStatusReg2[24]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[24]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[24]\);
    
    \MOSI_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \MOSI_obuf/U0/DOUT1\, Y => 
        \MOSI_obuf/U0/DOUT\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[30]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[30]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1061\, Y => 
        \MemorySynchronizer_0/N_1092\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_Y\, B
         => \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => ADLIB_GND0, S
         => OPEN, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0_Y\, 
        FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0_Z\, 
        CC => NET_CC_CONFIG627, P => NET_CC_CONFIG625, UB => 
        NET_CC_CONFIG626);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[8]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_8_S\, 
        Y => \MemorySynchronizer_0/N_2430\);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.un151_in_enablelto31_1\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/temp_1[25]\, B => 
        \MemorySynchronizer_0/temp_1[26]\, C => 
        \MemorySynchronizer_0/temp_1[27]\, D => 
        \MemorySynchronizer_0/temp_1[28]\, Y => 
        \MemorySynchronizer_0/un151_in_enablelto31_1\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_205\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_GND0, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1]\, 
        IPC => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WLAST_net\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_47_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[0]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_47\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[4]\, B => 
        \MemorySynchronizer_0/un104_in_enable_4\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[4]\);
    
    \STAMP_0/spi_dms2_cs\ : SLE
      port map(D => \STAMP_0/spi_dms2_cs_13_iv_i_Z\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/N_46\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => stamp0_spi_dms2_cs_c);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_144\ : 
        IP_INTERFACE
      port map(A => \sb_sb_0/FIC_0_LOCK\, B => ADLIB_VCC1, C => 
        ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_46_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_66\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_46_set_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[2]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[2]\, 
        B => \sb_sb_0_STAMP_PWDATA[2]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[2]\);
    
    \STAMP_0/delay_counter[4]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[4]\);
    
    \STAMP_0/un1_presetn_inv\ : CFG4
      generic map(INIT => x"FF7F")

      port map(A => \STAMP_0/un85_paddr_3_Z\, B => 
        debug_led_net_0, C => \STAMP_0/component_state_Z[3]\, D
         => sb_sb_0_STAMP_PWRITE, Y => 
        \STAMP_0/un1_presetn_inv_Z\);
    
    \STAMP_0/delay_counter_cry[8]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[8]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/delay_counter_cry_Z[7]\, S => 
        \STAMP_0/delay_counter_s[8]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[8]\, CC => NET_CC_CONFIG419, 
        P => NET_CC_CONFIG417, UB => NET_CC_CONFIG418);
    
    \STAMP_0/async_state_17_iv_0_RNO[1]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \STAMP_0/N_204\, B => 
        \STAMP_0/async_state_Z[0]\, Y => \STAMP_0/N_206\);
    
    \MemorySynchronizer_0/TimeStampGen/prescaler[4]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_5_Z[4]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[4]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[17]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[17]\, B => 
        \sb_sb_0_Memory_PRDATA[17]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[17]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[3]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[3]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1088\, Y => 
        \MemorySynchronizer_0/N_1119\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[3]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[3]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[2]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[3]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[3]\, CC
         => NET_CC_CONFIG15, P => NET_CC_CONFIG13, UB => 
        NET_CC_CONFIG14);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[21]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_21_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_88\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_139\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net\, IPB
         => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1]\, 
        IPC => OPEN);
    
    \STAMP_0/dummy[7]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_67\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[7]\);
    
    \RXSM_SODS_ibuf/U0/U_IOINFF\ : IOINFF_BYPASS
      port map(A => \RXSM_SODS_ibuf/U0/YIN1\, Y => 
        \RXSM_SODS_ibuf/U0/YIN\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_0_a1_Z\, 
        B => \MemorySynchronizer_0/N_140_2\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_4_Z\, 
        D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a0_1_Z\, 
        Y => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\);
    
    \debug_led_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \debug_led_obuf/U0/DOUT1\, Y => 
        \debug_led_obuf/U0/DOUT\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_7\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[7]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_6_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[7]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_7_Z\, 
        CC => NET_CC_CONFIG125, P => NET_CC_CONFIG123, UB => 
        NET_CC_CONFIG124);
    
    \STAMP_0/un1_component_state_9_i_o2_0\ : CFG2
      generic map(INIT => x"B")

      port map(A => \STAMP_0/spi_busy\, B => 
        \STAMP_0/component_state_Z[1]\, Y => \STAMP_0/N_160\);
    
    \STAMP_0/measurement_dms2[0]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[32]\);
    
    \STAMP_0/spi/count_cry[18]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[18]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[17]\, S => 
        \STAMP_0/spi/count_s[18]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[18]\, CC => NET_CC_CONFIG979, P
         => NET_CC_CONFIG977, UB => NET_CC_CONFIG978);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_135\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net\, 
        IPC => OPEN);
    
    \STAMP_0/un45_async_state_cry_4\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \STAMP_0/config_Z[28]\, B => 
        \STAMP_0_data_frame[7]\, C => ADLIB_GND0, D => ADLIB_GND0, 
        FCI => \STAMP_0/un45_async_state_cry_3_Z\, S => OPEN, Y
         => OPEN, FCO => \STAMP_0/un45_async_state_cry_4_Z\, CC
         => NET_CC_CONFIG528, P => NET_CC_CONFIG526, UB => 
        NET_CC_CONFIG527);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_23\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[23]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_22_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_23_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_23_Z\, 
        CC => NET_CC_CONFIG696, P => NET_CC_CONFIG694, UB => 
        NET_CC_CONFIG695);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[24]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[24]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[24]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[24]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[24]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[24]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[12]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[12]\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/N_2323\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[12]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[12]\);
    
    \STAMP_0/un1_spi_rx_data_0[25]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame[25]\, B => 
        \STAMP_0/config_Z[25]\, C => \sb_sb_0_STAMP_PADDR[8]\, Y
         => \STAMP_0/N_608\);
    
    \STAMP_0/delay_counter[26]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[26]\);
    
    \STAMP_0/un1_spi_rx_data_2[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_586\, B => \STAMP_0/N_620\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_653\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[14]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[14]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[14]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[14]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_0_a1_Z\, 
        B => \MemorySynchronizer_0/N_140_2\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_4_Z\, 
        D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a0_1_Z\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_Z\);
    
    \STAMP_0/spi/count[31]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[31]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB12_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[31]\);
    
    \stamp0_spi_dms2_cs_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \stamp0_spi_dms2_cs_obuf/U0/DOUT1\, Y => 
        \stamp0_spi_dms2_cs_obuf/U0/DOUT\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[8]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[8]\, 
        B => \sb_sb_0_STAMP_PWDATA[8]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[8]\);
    
    \MemorySynchronizer_0/waitingtimercounter_RNIA97L[26]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_46_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[26]\, C
         => \MemorySynchronizer_0/un1_nreset_39_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[26]\);
    
    \MemorySynchronizer_0/PRDATA[26]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[26]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[26]\);
    
    \MemorySynchronizer_0/un1_nreset_30\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[4]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_30_i\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[31]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2585\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[31]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[31]\, D => 
        \MemorySynchronizer_0/N_1201\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[31]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_9\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[9]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_8_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_9_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_9_Z\, CC
         => NET_CC_CONFIG752, P => NET_CC_CONFIG750, UB => 
        NET_CC_CONFIG751);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[31]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[31]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[31]\);
    
    \STAMP_0/new_avail_0_sqmuxa_1_0_a3\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \STAMP_0_data_frame[15]\, B => 
        \STAMP_0_data_frame[14]\, C => \STAMP_0/config_Z[30]\, D
         => \STAMP_0/N_333\, Y => \STAMP_0/new_avail_0_sqmuxa_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_o2[19]\ : CFG4
      generic map(INIT => x"F2F0")

      port map(A => \MemorySynchronizer_0/N_2316\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2572\, D => 
        \MemorySynchronizer_0/N_271\, Y => 
        \MemorySynchronizer_0/N_2323\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_150\ : 
        IP_INTERFACE
      port map(A => RXSM_SODS_c, B => MISO_c, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_RNI8TKQ[28]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_44_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[28]\, C
         => \MemorySynchronizer_0/un1_nreset_37_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[28]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[7]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_7\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[7]\, 
        C => \MemorySynchronizer_0/N_1545\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[7]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[4]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[4]\, B => 
        \sb_sb_0_STAMP_PWDATA[4]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[4]\);
    
    \STAMP_0/spi/tx_buffer_RNO[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[10]\, B => 
        \STAMP_0/spi/tx_buffer_Z[9]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_125\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[9]\ : SLE
      port map(D => \STAMP_0_data_frame[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[9]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_22\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[22]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_21_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[10]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_22_Z\, CC
         => NET_CC_CONFIG363, P => NET_CC_CONFIG361, UB => 
        NET_CC_CONFIG362);
    
    \MemorySynchronizer_0/TimeStampGen/counter[26]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[26]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[26]\);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB8\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\);
    
    \MemorySynchronizer_0/TimeStampReg[31]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[31]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[31]\);
    
    \MemorySynchronizer_0/waitingtimercounter[26]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[26]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_39_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[26]\);
    
    \MemorySynchronizer_0/un1_nreset_57_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_57_i_i_a2_Z\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_57_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_57_rs_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/prescaler[1]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc1_Z\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[1]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_6\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[6]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_5_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[26]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_6_Z\, CC
         => NET_CC_CONFIG315, P => NET_CC_CONFIG313, UB => 
        NET_CC_CONFIG314);
    
    \MemorySynchronizer_0/resynctimercounter[19]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1103\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[19]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_63\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[1]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[1]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_s_387_FCO\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[1]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[1]\, CC
         => NET_CC_CONFIG9, P => NET_CC_CONFIG7, UB => 
        NET_CC_CONFIG8);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_8\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[8]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[8]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_7\, S => 
        \MemorySynchronizer_0/temp_1[8]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_8\, CC => 
        NET_CC_CONFIG223, P => NET_CC_CONFIG221, UB => 
        NET_CC_CONFIG222);
    
    AFLSDF_INV_5 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_5\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[12]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[12]\, B => 
        \sb_sb_0_Memory_PRDATA[12]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12]\);
    
    \ResetAND_RNIMHJB/U0_RGB1\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_YR\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_136\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net\, IPB
         => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un104_in_enable_cry_0_CC_0\ : CC_CONFIG
      port map(CI => ADLIB_GND0, CO => CI_TO_CO819, P(0) => 
        NET_CC_CONFIG821, P(1) => NET_CC_CONFIG824, P(2) => 
        NET_CC_CONFIG827, P(3) => NET_CC_CONFIG830, P(4) => 
        NET_CC_CONFIG833, P(5) => NET_CC_CONFIG836, P(6) => 
        NET_CC_CONFIG839, P(7) => NET_CC_CONFIG842, P(8) => 
        NET_CC_CONFIG845, P(9) => NET_CC_CONFIG848, P(10) => 
        NET_CC_CONFIG851, P(11) => NET_CC_CONFIG854, UB(0) => 
        NET_CC_CONFIG822, UB(1) => NET_CC_CONFIG825, UB(2) => 
        NET_CC_CONFIG828, UB(3) => NET_CC_CONFIG831, UB(4) => 
        NET_CC_CONFIG834, UB(5) => NET_CC_CONFIG837, UB(6) => 
        NET_CC_CONFIG840, UB(7) => NET_CC_CONFIG843, UB(8) => 
        NET_CC_CONFIG846, UB(9) => NET_CC_CONFIG849, UB(10) => 
        NET_CC_CONFIG852, UB(11) => NET_CC_CONFIG855, CC(0) => 
        NET_CC_CONFIG823, CC(1) => NET_CC_CONFIG826, CC(2) => 
        NET_CC_CONFIG829, CC(3) => NET_CC_CONFIG832, CC(4) => 
        NET_CC_CONFIG835, CC(5) => NET_CC_CONFIG838, CC(6) => 
        NET_CC_CONFIG841, CC(7) => NET_CC_CONFIG844, CC(8) => 
        NET_CC_CONFIG847, CC(9) => NET_CC_CONFIG850, CC(10) => 
        NET_CC_CONFIG853, CC(11) => NET_CC_CONFIG856);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[26]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_26\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[26]\, 
        C => \MemorySynchronizer_0/N_1493\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[26]\);
    
    \MemorySynchronizer_0/un1_nreset_51_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_38\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_51_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_51_rs_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[19]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[19]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[19]\);
    
    \STAMP_0/un1_presetn_inv_RNIK8BR\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/un1_presetn_inv_Z\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_5\, Y => 
        \STAMP_0/un1_presetn_inv_RNIK8BR_Z\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_8\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/PWRITE_net\, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX2_SEL_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[6]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_234\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg[2]\ : SLE
      port map(D => \MemorySynchronizer_0/SynchStatusReg_168[0]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, 
        EN => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[2]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[6]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[6]\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_6_S\, 
        C => \MemorySynchronizer_0/resettimercounter_m[6]\, D => 
        \MemorySynchronizer_0/resettimercounter_0_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9[6]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[26]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[26]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1065\, Y => 
        \MemorySynchronizer_0/N_1096\);
    
    \STAMP_0/measurement_dms1[0]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[48]\);
    
    AFLSDF_INV_64 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_43_Z\, Y => 
        \AFLSDF_INV_64\);
    
    \STAMP_0/un1_spi_rx_data_1[8]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[40]\, B => 
        \STAMP_0/dummy_Z[8]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_625\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_24\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[24]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_23_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[8]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_24_Z\, CC
         => NET_CC_CONFIG369, P => NET_CC_CONFIG367, UB => 
        NET_CC_CONFIG368);
    
    \MemorySynchronizer_0/un1_nreset_24_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_61\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_24_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_24_rs_Z\);
    
    \STAMP_0/un1_spi_rx_data_1[28]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[60]\, B => 
        \STAMP_0/dummy_Z[28]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_645\);
    
    \STAMP_0/un1_spi_rx_data_1[12]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[44]\, B => 
        \STAMP_0/dummy_Z[12]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_629\);
    
    \STAMP_0/async_prescaler_count_5[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/un1_async_prescaler_count\, B => 
        \STAMP_0/un5_async_prescaler_count_s_11_S\, Y => 
        \STAMP_0/async_prescaler_count_5_Z[11]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[19]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_19\);
    
    \STAMP_0/delay_counter_cry[1]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[1]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/delay_counter_cry_Z[0]\, S => 
        \STAMP_0/delay_counter_s[1]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[1]\, CC => NET_CC_CONFIG398, 
        P => NET_CC_CONFIG396, UB => NET_CC_CONFIG397);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[20]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[20]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[12]\, Y
         => \MemorySynchronizer_0/N_1071\);
    
    \STAMP_0/status_dms1_overwrittenVal_RNO\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/un1_new_avail_0_sqmuxa_1\, B => 
        \STAMP_0_data_frame[15]\, Y => \STAMP_0/N_116_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_10\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15]\, C
         => ADLIB_VCC1, IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15]\, 
        IPC => OPEN);
    
    \STAMP_0/spi/mosi_cl\ : SLE
      port map(D => \STAMP_0/spi/N_25_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => mosi_cl);
    
    \STAMP_0/config[8]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[8]\);
    
    \STAMP_0/un1_component_state_13_i_0\ : CFG4
      generic map(INIT => x"D000")

      port map(A => \STAMP_0/component_state_Z[0]\, B => 
        \STAMP_0/un1_component_state_13_i_a3_0_0_Z\, C => 
        \STAMP_0/N_164\, D => \STAMP_0/N_337\, Y => 
        \STAMP_0/un1_component_state_13_i_0_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_o2[10]\ : CFG4
      generic map(INIT => x"1FF8")

      port map(A => \sb_sb_0_STAMP_PADDR[2]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, C => \sb_sb_0_STAMP_PADDR[4]\, 
        D => \sb_sb_0_STAMP_PADDR[5]\, Y => 
        \MemorySynchronizer_0/N_2317\);
    
    \STAMP_0/status_async_cycles[1]\ : SLE
      port map(D => \STAMP_0/status_async_cycles_lm[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/status_async_cycles_1_sqmuxa_1_i_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[4]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[3]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[3]\);
    
    \STAMP_0/delay_counter[19]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[19]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS_1[0]\ : CFG4
      generic map(INIT => x"7000")

      port map(A => \sb_sb_0/STAMP_PADDRS[14]\, B => 
        \sb_sb_0/STAMP_PADDRS[13]\, C => 
        \sb_sb_0/CoreAPB3_0/iPSELS_raw_1_0_Z[0]\, D => 
        \sb_sb_0/STAMP_PADDRS[12]\, Y => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS[0]\);
    
    \MemorySynchronizer_0/TimeStampReg[29]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[29]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[29]\);
    
    \STAMP_0/measurement_temp[3]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[19]\);
    
    \STAMP_0/spi/rx_buffer_0_sqmuxa_1_0_o2\ : CFG4
      generic map(INIT => x"7555")

      port map(A => \STAMP_0/spi/clk_toggles_Z[5]\, B => 
        \STAMP_0/spi/clk_toggles_Z[0]\, C => 
        \STAMP_0/spi/un10_count_0_a2_0_Z\, D => 
        \STAMP_0/spi/un10_count_0_a2_0_0_Z\, Y => 
        \STAMP_0/spi/N_30\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[0]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[0]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1091\, Y => 
        \MemorySynchronizer_0/N_1122\);
    
    \adc_clk_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => adc_clk, D => \adc_clk_obuf/U0/DOUT\, E => 
        \adc_clk_obuf/U0/EOUT\);
    
    \STAMP_0/un1_spi_rx_data_2[21]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_604\, B => \STAMP_0/N_638\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_671\);
    
    \MemorySynchronizer_0/ResetTimerValueReg_RNIJ7VC[11]\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[11]\, B => 
        NN_1, Y => \MemorySynchronizer_0/N_21_i\);
    
    \STAMP_0/un85_paddr_3\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \STAMP_0/un52_paddr_2_1\, B => 
        \STAMP_0/un76_paddr_0_a2_2_Z\, C => 
        \STAMP_0/un52_paddr_2_0_Z\, D => 
        \STAMP_0/un85_paddr_3_0_tz_Z\, Y => 
        \STAMP_0/un85_paddr_3_Z\);
    
    AFLSDF_INV_73 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_35_Z\, Y => 
        \AFLSDF_INV_73\);
    
    \STAMP_0/spi/un7_count_NE_23\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \STAMP_0/spi/count_Z[23]\, B => 
        \STAMP_0/spi/count_Z[22]\, C => \STAMP_0/spi/count_Z[21]\, 
        D => \STAMP_0/spi/count_Z[20]\, Y => 
        \STAMP_0/spi/un7_count_NE_23_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[15]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[15]\, B => 
        \sb_sb_0_STAMP_PWDATA[15]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[15]\);
    
    \MemorySynchronizer_0/PRDATA[2]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[2]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[2]\);
    
    \STAMP_0/PRDATA[13]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[13]\);
    
    \STAMP_0/un5_async_prescaler_count_cry_6\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[6]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_5_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_6_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_6_Z\, CC
         => NET_CC_CONFIG498, P => NET_CC_CONFIG496, UB => 
        NET_CC_CONFIG497);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_51_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[25]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_51\);
    
    \MemorySynchronizer_0/SynchStatusReg2[30]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[30]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[30]\);
    
    \STAMP_0/async_state_RNO[0]\ : CFG4
      generic map(INIT => x"0041")

      port map(A => \STAMP_0/un1_async_state_0_sqmuxa_i\, B => 
        \STAMP_0/N_204\, C => \STAMP_0/async_state_Z[0]\, D => 
        \STAMP_0/request_resync_1_sqmuxa_1_Z\, Y => 
        \STAMP_0/N_90_i\);
    
    \MemorySynchronizer_0/TimeStampReg[4]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[4]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[4]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[23]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_84\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[23]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[23]\, 
        D => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[23]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_12\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_13\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_11_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[13]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_12_Z\, CC
         => NET_CC_CONFIG1059, P => NET_CC_CONFIG1057, UB => 
        NET_CC_CONFIG1058);
    
    \MemorySynchronizer_0/resynceventpulldowncounter[0]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1158_i_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[0]\);
    
    \stamp0_spi_dms2_cs_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => stamp0_spi_dms2_cs, D => 
        \stamp0_spi_dms2_cs_obuf/U0/DOUT\, E => 
        \stamp0_spi_dms2_cs_obuf/U0/EOUT\);
    
    \STAMP_0/measurement_temp[2]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[18]\);
    
    \STAMP_0/delay_counter_RNIG01L3[16]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \STAMP_0/N_517_i_0_a2_14\, B => 
        \STAMP_0/N_517_i_0_a2_25\, C => \STAMP_0/N_517_i_0_a2_20\, 
        D => \STAMP_0/N_517_i_0_a2_15\, Y => \STAMP_0/N_238\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_0_CC_2\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO722, CO => OPEN, P(0) => 
        NET_CC_CONFIG795, P(1) => NET_CC_CONFIG798, P(2) => 
        NET_CC_CONFIG801, P(3) => NET_CC_CONFIG804, P(4) => 
        NET_CC_CONFIG807, P(5) => NET_CC_CONFIG810, P(6) => 
        NET_CC_CONFIG813, P(7) => NET_CC_CONFIG816, P(8) => 
        ADLIB_VCC1, P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, 
        P(11) => ADLIB_VCC1, UB(0) => NET_CC_CONFIG796, UB(1) => 
        NET_CC_CONFIG799, UB(2) => NET_CC_CONFIG802, UB(3) => 
        NET_CC_CONFIG805, UB(4) => NET_CC_CONFIG808, UB(5) => 
        NET_CC_CONFIG811, UB(6) => NET_CC_CONFIG814, UB(7) => 
        NET_CC_CONFIG817, UB(8) => ADLIB_VCC1, UB(9) => 
        ADLIB_VCC1, UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, 
        CC(0) => NET_CC_CONFIG797, CC(1) => NET_CC_CONFIG800, 
        CC(2) => NET_CC_CONFIG803, CC(3) => NET_CC_CONFIG806, 
        CC(4) => NET_CC_CONFIG809, CC(5) => NET_CC_CONFIG812, 
        CC(6) => NET_CC_CONFIG815, CC(7) => NET_CC_CONFIG818, 
        CC(8) => nc332, CC(9) => nc81, CC(10) => nc375, CC(11)
         => nc201);
    
    \STAMP_0/async_state_1_sqmuxa_i_o3_RNINQM71\ : CFG4
      generic map(INIT => x"FEFF")

      port map(A => \STAMP_0/component_state_Z[1]\, B => 
        \STAMP_0/component_state_Z[5]\, C => \STAMP_0/N_163\, D
         => \STAMP_0/N_197\, Y => \STAMP_0/N_204\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_11[28]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \sb_sb_0_STAMP_PADDR[5]\, B => 
        \MemorySynchronizer_0/N_2575\, C => 
        \sb_sb_0_STAMP_PADDR[4]\, Y => 
        \MemorySynchronizer_0/N_2593\);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_27\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_17_Z\, B => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_16_Z\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_15_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_18_Z\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_36\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[5]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[7]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[5]\, C => 
        \MemorySynchronizer_0/N_2576\, D => 
        \MemorySynchronizer_0/N_1182\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[5]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[26]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[26]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[26]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[26]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[26]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[26]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[28]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[28]\);
    
    \STAMP_0/un1_spi_rx_data_1[4]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[36]\, B => 
        \STAMP_0/dummy_Z[4]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_621\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_101\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[1]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[8]\, 
        IPC => OPEN);
    
    \STAMP_0/spi/clk_toggles[0]\ : SLE
      port map(D => \STAMP_0/spi/clk_toggles_lm[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB14_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_37_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/clk_toggles_Z[0]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[21]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[21]\, B => 
        \sb_sb_0_STAMP_PWDATA[21]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[21]\);
    
    AFLSDF_INV_76 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_76\);
    
    \STAMP_0/async_prescaler_count_5[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \STAMP_0/un1_async_prescaler_count\, B => 
        \STAMP_0/async_prescaler_count_Z[0]\, Y => 
        \STAMP_0/async_prescaler_count_5_Z[0]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[1]\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[1]\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[1]\, C => 
        \MemorySynchronizer_0/N_2593\, D => 
        \MemorySynchronizer_0/N_1172\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[1]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_0_CC_0\ : 
        CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => CI_TO_CO1019, P(0) => 
        ADLIB_VCC1, P(1) => ADLIB_VCC1, P(2) => ADLIB_GND0, P(3)
         => NET_CC_CONFIG1021, P(4) => NET_CC_CONFIG1024, P(5)
         => NET_CC_CONFIG1027, P(6) => NET_CC_CONFIG1030, P(7)
         => NET_CC_CONFIG1033, P(8) => NET_CC_CONFIG1036, P(9)
         => NET_CC_CONFIG1039, P(10) => NET_CC_CONFIG1042, P(11)
         => NET_CC_CONFIG1045, UB(0) => ADLIB_VCC1, UB(1) => 
        ADLIB_VCC1, UB(2) => ADLIB_VCC1, UB(3) => 
        NET_CC_CONFIG1022, UB(4) => NET_CC_CONFIG1025, UB(5) => 
        NET_CC_CONFIG1028, UB(6) => NET_CC_CONFIG1031, UB(7) => 
        NET_CC_CONFIG1034, UB(8) => NET_CC_CONFIG1037, UB(9) => 
        NET_CC_CONFIG1040, UB(10) => NET_CC_CONFIG1043, UB(11)
         => NET_CC_CONFIG1046, CC(0) => nc168, CC(1) => nc425, 
        CC(2) => nc323, CC(3) => NET_CC_CONFIG1023, CC(4) => 
        NET_CC_CONFIG1026, CC(5) => NET_CC_CONFIG1029, CC(6) => 
        NET_CC_CONFIG1032, CC(7) => NET_CC_CONFIG1035, CC(8) => 
        NET_CC_CONFIG1038, CC(9) => NET_CC_CONFIG1041, CC(10) => 
        NET_CC_CONFIG1044, CC(11) => NET_CC_CONFIG1047);
    
    \MemorySynchronizer_0/waitingtimercounter[30]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[30]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_35_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[30]\);
    
    \MemorySynchronizer_0/TimeStampReg[19]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[19]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[19]\);
    
    \MemorySynchronizer_0/ConfigReg[22]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[22]\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_213\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1]\, 
        IPC => OPEN);
    
    AND2_0 : CFG2
      generic map(INIT => x"8")

      port map(A => NN_1, B => ADLIB_VCC1, Y => debug_led_net_0);
    
    \STAMP_0/un76_paddr_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/un76_paddr_0_a2_2_Z\, B => 
        \STAMP_0/un52_paddr_2_0_Z\, Y => \STAMP_0/un76_paddr\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_20\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[25]\, B
         => ADLIB_GND0, C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net\, 
        IPC => OPEN);
    
    AFLSDF_INV_28 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_28\);
    
    \STAMP_0/async_prescaler_count[9]\ : SLE
      port map(D => \STAMP_0/un5_async_prescaler_count_cry_9_S\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[9]\);
    
    AFLSDF_INV_88 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_57_i_i_a2_Z\, 
        Y => \AFLSDF_INV_88\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_s_31\ : 
        ARI1_CC
      generic map(INIT => x"49900")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_axb_31\, C => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, D
         => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_30_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_s_31_S\, 
        Y => OPEN, FCO => OPEN, CC => NET_CC_CONFIG720, P => 
        NET_CC_CONFIG718, UB => NET_CC_CONFIG719);
    
    \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa_i_0_i_a2\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa_i_0_i_a2_1_Z\, 
        B => \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[4]\, D => \sb_sb_0_STAMP_PADDR[5]\, 
        Y => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\);
    
    \MemorySynchronizer_0/un1_nreset_59_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[7]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_59_i\);
    
    \STAMP_0/un1_spi_rx_data_0[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[6]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[6]\, Y
         => \STAMP_0/N_589\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[19]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_19_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[13]\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO[27]\ : CFG4
      generic map(INIT => x"0F0B")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[27]\, 
        B => \MemorySynchronizer_0/MemorySyncState_Z[3]\, C => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_0_a2_0_0_Z[25]\, 
        D => \MemorySynchronizer_0/N_2321\, Y => 
        \MemorySynchronizer_0/N_2035_i\);
    
    \MemorySynchronizer_0/SynchStatusReg2[7]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[7]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[7]\);
    
    \MemorySynchronizer_0/un1_nreset_19_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_32_i_i_a2_Z\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_19_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_19_rs_Z\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_28\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_19_Z\, 
        B => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_16_Z\, 
        C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_17_Z\, 
        D => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_18_Z\, 
        Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_28_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_230\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter[19]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_14_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[19]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_21\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_22\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_20_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[22]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_21_Z\, CC
         => NET_CC_CONFIG1086, P => NET_CC_CONFIG1084, UB => 
        NET_CC_CONFIG1085);
    
    \adc_start_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \adc_start_obuf/U0/EOUT1\, Y => 
        \adc_start_obuf/U0/EOUT\);
    
    \STAMP_0/un76_paddr_0_a2_2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \sb_sb_0_STAMP_PADDR[9]\, B => 
        \sb_sb_0_STAMP_PADDR[7]\, C => \STAMP_0/un52_paddr_2_Z\, 
        D => \STAMP_0/un52_paddr_5_Z\, Y => 
        \STAMP_0/un76_paddr_0_a2_2_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_112\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1]\, 
        IPC => OPEN);
    
    \STAMP_0/delay_counter_lm_0[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[8]\, Y => 
        \STAMP_0/delay_counter_lm[8]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[1]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[1]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[1]\, D => 
        \MemorySynchronizer_0/un5_resettimercounter_m[31]\, Y => 
        \MemorySynchronizer_0/resettimercounter_9[1]\);
    
    \STAMP_0/measurement_dms1[6]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[54]\);
    
    \STAMP_0/un1_component_state_9_i_o2\ : CFG3
      generic map(INIT => x"73")

      port map(A => \STAMP_0/apb_spi_finished_Z\, B => 
        \STAMP_0/component_state_Z[3]\, C => 
        \STAMP_0/un13_paddr_i_0\, Y => \STAMP_0/N_155\);
    
    \STAMP_0/config[9]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[9]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[9]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[9]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[9]\, C => 
        \MemorySynchronizer_0/N_2576\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[9]\);
    
    \STAMP_0/un1_spi_rx_data_1[6]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[38]\, B => 
        \STAMP_0/dummy_Z[6]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_623\);
    
    \STAMP_0/spi/clk_toggles_s[5]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/spi/clk_toggles_Z[5]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/spi/clk_toggles_cry_Z[4]\, S
         => \STAMP_0/spi/clk_toggles_s_Z[5]\, Y => OPEN, FCO => 
        OPEN, CC => NET_CC_CONFIG622, P => NET_CC_CONFIG620, UB
         => NET_CC_CONFIG621);
    
    \MemorySynchronizer_0/un1_nreset_40_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[19]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_40_i\);
    
    \adc_clk_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \adc_clk_obuf/U0/DOUT1\, Y => 
        \adc_clk_obuf/U0/DOUT\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[27]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[27]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[27]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[5]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[27]\);
    
    \MemorySynchronizer_0/resettimercounter[2]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[2]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_32_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[2]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv[5]\ : CFG4
      generic map(INIT => x"FBFA")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_m[7]\, B
         => STAMP_0_new_avail, C => 
        \MemorySynchronizer_0/SynchStatusReg_82_m[5]\, D => 
        \MemorySynchronizer_0/N_1512\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168[5]\);
    
    \STAMP_0/config[16]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[16]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[5]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[5]\, B => 
        \sb_sb_0_Memory_PRDATA[5]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5]\);
    
    \MemorySynchronizer_0/ConfigReg[3]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[3]\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_57\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[19]\, B => 
        \MemorySynchronizer_0/un104_in_enable_18\, C => 
        \MemorySynchronizer_0/un104_in_enable_19\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[18]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[8]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[9]\, CC
         => NET_CC_CONFIG565, P => NET_CC_CONFIG563, UB => 
        NET_CC_CONFIG564);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0[30]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/N_1222\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[30]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[30]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[30]\, Y => 
        \MemorySynchronizer_0/PRDATA_21[30]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[26]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[26]\, B => 
        \sb_sb_0_Memory_PRDATA[26]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[26]\);
    
    \MemorySynchronizer_0/PRDATA[10]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[10]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[10]\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0[1]\ : CFG4
      generic map(INIT => x"BAAA")

      port map(A => 
        \MemorySynchronizer_0/MemorySyncState_ns_0_0_Z[1]\, B => 
        STAMP_0_new_avail, C => 
        \MemorySynchronizer_0/un41_in_enable_i_0\, D => 
        \MemorySynchronizer_0/N_1495\, Y => 
        \MemorySynchronizer_0/MemorySyncState_ns[1]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_22\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[22]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[22]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_21_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_22_Z\, CC => 
        NET_CC_CONFIG889, P => NET_CC_CONFIG887, UB => 
        NET_CC_CONFIG888);
    
    \MemorySynchronizer_0/TimeStampGen/counter[22]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[22]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[22]\);
    
    \STAMP_0/delay_counter_cry[0]_CC_1\ : CC_CONFIG
      port map(CI => CI_TO_CO391, CO => CI_TO_CO392, P(0) => 
        NET_CC_CONFIG429, P(1) => NET_CC_CONFIG432, P(2) => 
        NET_CC_CONFIG435, P(3) => NET_CC_CONFIG438, P(4) => 
        NET_CC_CONFIG441, P(5) => NET_CC_CONFIG444, P(6) => 
        NET_CC_CONFIG447, P(7) => NET_CC_CONFIG450, P(8) => 
        NET_CC_CONFIG453, P(9) => NET_CC_CONFIG456, P(10) => 
        NET_CC_CONFIG459, P(11) => NET_CC_CONFIG462, UB(0) => 
        NET_CC_CONFIG430, UB(1) => NET_CC_CONFIG433, UB(2) => 
        NET_CC_CONFIG436, UB(3) => NET_CC_CONFIG439, UB(4) => 
        NET_CC_CONFIG442, UB(5) => NET_CC_CONFIG445, UB(6) => 
        NET_CC_CONFIG448, UB(7) => NET_CC_CONFIG451, UB(8) => 
        NET_CC_CONFIG454, UB(9) => NET_CC_CONFIG457, UB(10) => 
        NET_CC_CONFIG460, UB(11) => NET_CC_CONFIG463, CC(0) => 
        NET_CC_CONFIG431, CC(1) => NET_CC_CONFIG434, CC(2) => 
        NET_CC_CONFIG437, CC(3) => NET_CC_CONFIG440, CC(4) => 
        NET_CC_CONFIG443, CC(5) => NET_CC_CONFIG446, CC(6) => 
        NET_CC_CONFIG449, CC(7) => NET_CC_CONFIG452, CC(8) => 
        NET_CC_CONFIG455, CC(9) => NET_CC_CONFIG458, CC(10) => 
        NET_CC_CONFIG461, CC(11) => NET_CC_CONFIG464);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_2\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[2]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[2]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_1\, S => 
        \MemorySynchronizer_0/temp_1[2]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_2\, CC => 
        NET_CC_CONFIG205, P => NET_CC_CONFIG203, UB => 
        NET_CC_CONFIG204);
    
    \stamp0_ready_dms2_ibuf/U0/U_IOINFF\ : IOINFF_BYPASS
      port map(A => \stamp0_ready_dms2_ibuf/U0/YIN1\, Y => 
        \stamp0_ready_dms2_ibuf/U0/YIN\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_215\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3]\, 
        IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data[5]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_655\, C => \STAMP_0/spi_rx_data[5]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[5]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[4]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[4]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1[28]\, Y => 
        \MemorySynchronizer_0/N_1087\);
    
    \STAMP_0/delay_counter_cry[17]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[17]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[16]\, S
         => \STAMP_0/delay_counter_s[17]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[17]\, CC => NET_CC_CONFIG446, 
        P => NET_CC_CONFIG444, UB => NET_CC_CONFIG445);
    
    \MemorySynchronizer_0/un1_nreset_19_rs_RNIE5UN\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_2539_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[28]\, C => 
        \MemorySynchronizer_0/un1_nreset_19_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[28]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_45_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[27]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_45\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_209\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/MemorySyncState_RNIJVOS[3]\ : CFG3
      generic map(INIT => x"13")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => \MemorySynchronizer_0/un1_enabletimestampgen2_2_sn\, 
        C => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, Y
         => \MemorySynchronizer_0/N_2304_i\);
    
    \STAMP_0/config[28]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[28]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_15\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[15]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_14_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[15]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_15_Z\, 
        CC => NET_CC_CONFIG149, P => NET_CC_CONFIG147, UB => 
        NET_CC_CONFIG148);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[24]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_24\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[7]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[7]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[6]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[7]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[7]\, CC
         => NET_CC_CONFIG27, P => NET_CC_CONFIG25, UB => 
        NET_CC_CONFIG26);
    
    \MemorySynchronizer_0/ConfigReg[23]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[23]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[22]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[22]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[22]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[22]\);
    
    \STAMP_0/async_state_0_sqmuxa\ : CFG4
      generic map(INIT => x"0800")

      port map(A => MemorySynchronizer_0_dataReadyReset, B => 
        \STAMP_0/async_state_Z[0]\, C => 
        \STAMP_0/async_state_Z[1]\, D => 
        \STAMP_0/component_state_Z[5]\, Y => 
        \STAMP_0/async_state_0_sqmuxa_Z\);
    
    \MemorySynchronizer_0/SynchronizerInterrupt\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa_i\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, 
        EN => 
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa_1_i_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        MemorySynchronizer_0_SynchronizerInterrupt);
    
    \MemorySynchronizer_0/ConfigReg[19]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[19]\);
    
    \STAMP_0/measurement_dms1[1]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[49]\);
    
    \STAMP_0/spi/count_cry[20]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[20]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[19]\, S => 
        \STAMP_0/spi/count_s[20]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[20]\, CC => NET_CC_CONFIG985, P
         => NET_CC_CONFIG983, UB => NET_CC_CONFIG984);
    
    \MemorySynchronizer_0/SynchStatusReg2[12]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[12]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[12]\);
    
    \STAMP_0/measurement_temp[12]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[28]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_26\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[26]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[26]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_25\, S => 
        \MemorySynchronizer_0/temp_1[26]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_26\, CC => 
        NET_CC_CONFIG277, P => NET_CC_CONFIG275, UB => 
        NET_CC_CONFIG276);
    
    \MemorySynchronizer_0/un1_nreset_29_rs_RNI9THR\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_48_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[25]\, C => 
        \MemorySynchronizer_0/un1_nreset_29_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[25]\);
    
    \STAMP_0/dummy[23]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_68\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[23]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[2]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[2]\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0_o3_i_a2[1]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[2]\, B
         => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[1]\, C
         => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[0]\, Y
         => \MemorySynchronizer_0/N_2553\);
    
    \STAMP_0/un13_paddr\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \sb_sb_0_STAMP_PADDR[5]\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => sb_sb_0_STAMP_PWRITE, D
         => \sb_sb_0_STAMP_PADDR[4]\, Y => 
        \STAMP_0/un13_paddr_i_0\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[22]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[22]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[21]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[22]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[22]\, CC
         => NET_CC_CONFIG72, P => NET_CC_CONFIG70, UB => 
        NET_CC_CONFIG71);
    
    \MemorySynchronizer_0/un1_nreset_39_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_46\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_39_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_39_rs_Z\);
    
    \MemorySynchronizer_0/un1_nreset_20_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[0]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_20_i\);
    
    \STAMP_0/config[31]\ : SLE
      port map(D => \STAMP_0/config_8[31]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_component_state_6_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[31]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_51_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_69\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_51_set_Z\);
    
    \adc_start_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => adc_start, D => \adc_start_obuf/U0/DOUT\, E
         => \adc_start_obuf/U0/EOUT\);
    
    \STAMP_0/un1_spi_rx_data_0[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[4]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[4]\, Y
         => \STAMP_0/N_587\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_87\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[3]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_17\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[17]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_16_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[17]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_17_Z\, 
        CC => NET_CC_CONFIG155, P => NET_CC_CONFIG153, UB => 
        NET_CC_CONFIG154);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[26]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[26]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[26]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[6]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[26]\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[18]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[18]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1073\, Y => 
        \MemorySynchronizer_0/N_1104\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_59_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[7]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_59\);
    
    
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1_0_a2_RNIU0KO2\ : 
        CFG4
      generic map(INIT => x"5504")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, B => 
        \MemorySynchronizer_0/N_140_2\, C => 
        \MemorySynchronizer_0/numberofnewavails_RNIEAMF1_Z[0]\, D
         => \MemorySynchronizer_0/g2_0_0\, Y => 
        \MemorySynchronizer_0/N_2606\);
    
    \STAMP_0/un1_spi_rx_data_2[7]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_590\, B => \STAMP_0/N_624\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_657\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[22]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[22]\, B => 
        \sb_sb_0_STAMP_PWDATA[22]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[22]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_6\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_7\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_5_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[7]\, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_6_Z\, 
        CC => NET_CC_CONFIG1041, P => NET_CC_CONFIG1039, UB => 
        NET_CC_CONFIG1040);
    
    \STAMP_0/delay_counter[1]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[1]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_19[20]\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[21]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[19]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[11]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[3]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_19_Z[20]\);
    
    \MemorySynchronizer_0/TimeStampReg[20]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[20]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[20]\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO[29]\ : CFG3
      generic map(INIT => x"32")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[29]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, C
         => \MemorySynchronizer_0/N_122_i\, Y => 
        \MemorySynchronizer_0/N_113_i\);
    
    \stamp0_spi_mosi_obuft/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => stamp0_spi_mosi, D => 
        \stamp0_spi_mosi_obuft/U0/DOUT\, E => 
        \stamp0_spi_mosi_obuft/U0/EOUT\);
    
    \STAMP_0/spi/clk_toggles[4]\ : SLE
      port map(D => \STAMP_0/spi/clk_toggles_lm[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB14_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_37_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/clk_toggles_Z[4]\);
    
    \STAMP_0/delay_counter_lm_0[14]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[14]\, Y => 
        \STAMP_0/delay_counter_lm[14]\);
    
    \STAMP_0/delay_counter[24]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[24]\);
    
    \STAMP_0/spi/count[11]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[11]\);
    
    \STAMP_0/delay_counter_cry[9]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[9]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/delay_counter_cry_Z[8]\, S => 
        \STAMP_0/delay_counter_s[9]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[9]\, CC => NET_CC_CONFIG422, 
        P => NET_CC_CONFIG420, UB => NET_CC_CONFIG421);
    
    \STAMP_0/un1_spi_rx_data_0[11]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[11]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[11]\, Y
         => \STAMP_0/N_594\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[19]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[19]\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2564\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1342\);
    
    \MemorySynchronizer_0/waitingtimercounter[10]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[10]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_56_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[10]\);
    
    \STAMP_0/spi/count[15]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[15]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_8\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[8]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_7_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[8]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_8_Z\, 
        CC => NET_CC_CONFIG128, P => NET_CC_CONFIG126, UB => 
        NET_CC_CONFIG127);
    
    \STAMP_0/spi/rx_data[3]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB0_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[3]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[3]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[3]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[5]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[3]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_40\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30]\, 
        IPC => OPEN);
    
    \STAMP_0/spi/ss_n_buffer_1_sqmuxa_0_a2\ : CFG3
      generic map(INIT => x"B3")

      port map(A => \STAMP_0/spi/un7_count_NE_i\, B => 
        \STAMP_0/spi/state_Z[0]\, C => \STAMP_0/spi/un10_count_i\, 
        Y => \STAMP_0/spi/ss_n_buffer_1_sqmuxa\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[29]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[29]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[29]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[3]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[29]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[3]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[3]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[3]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[3]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[20]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_20_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[12]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[16]\ : SLE
      port map(D => \STAMP_0_data_frame[48]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[16]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[30]\, B => 
        \sb_sb_0_STAMP_PWDATA[30]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[30]\);
    
    AFLSDF_INV_68 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_68\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[14]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[14]\, B => 
        \sb_sb_0_STAMP_PWDATA[14]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[14]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_11\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[16]\, C
         => ADLIB_VCC1, IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_194\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a1_0_0\ : 
        CFG3
      generic map(INIT => x"20")

      port map(A => \MemorySynchronizer_0/APBState_Z[0]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, C => \sb_sb_0_STAMP_PADDR[6]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a1_0_0_Z\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[5]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_5\);
    
    \STAMP_0/measurement_temp[13]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[29]\);
    
    \STAMP_0/status_async_cycles_lm_0[0]\ : CFG4
      generic map(INIT => x"0FEE")

      port map(A => \STAMP_0/status_async_cycles_2_sqmuxa\, B => 
        \STAMP_0/status_async_cycles_3_sqmuxa\, C => 
        \STAMP_0_data_frame[3]\, D => 
        \STAMP_0/status_async_cycles_1_sqmuxa_Z\, Y => 
        \STAMP_0/status_async_cycles_lm[0]\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_18\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_8_S\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_9_S\, 
        C => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_10_S\, D
         => \MemorySynchronizer_0/un5_resettimercounter_cry_11_S\, 
        Y => \MemorySynchronizer_0/un6_in_enable_0_a3_18_Z\);
    
    \STAMP_0/spi/tx_buffer[5]\ : SLE
      port map(D => \STAMP_0/spi/N_132\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[5]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[14]\ : SLE
      port map(D => \STAMP_0_data_frame[46]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[14]\);
    
    \STAMP_0/dummy[6]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_70\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[6]\);
    
    \MemorySynchronizer_0/resynctimercounter[0]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1122\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[0]\);
    
    \MemorySynchronizer_0/TimeStampReg[10]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[10]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[10]\);
    
    \MemorySynchronizer_0/un1_nreset_34_0_a3_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[0]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_34_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_237\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_24\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_25\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_23_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[25]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_24_Z\, CC
         => NET_CC_CONFIG1095, P => NET_CC_CONFIG1093, UB => 
        NET_CC_CONFIG1094);
    
    \MemorySynchronizer_0/ConfigReg[11]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[11]\);
    
    \MemorySynchronizer_0/un1_nreset_44_0_a3_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[9]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_44_i\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[24]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[3]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[24]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[24]\);
    
    \STAMP_0/spi_dms2_cs_1_sqmuxa_1_0_a3\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \STAMP_0/drdy_flank_detected_dms2_Z\, B => 
        \STAMP_0/drdy_flank_detected_dms1_Z\, C => 
        \STAMP_0/config_Z[30]\, D => \STAMP_0/N_333\, Y => 
        \STAMP_0/spi_dms2_cs_1_sqmuxa_1\);
    
    \MemorySynchronizer_0/SynchStatusReg[7]\ : SLE
      port map(D => \MemorySynchronizer_0/SynchStatusReg_168[5]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, 
        EN => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[7]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg_RNIK8VC[12]\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[12]\, B => 
        NN_1, Y => \MemorySynchronizer_0/N_1981_i\);
    
    \AND2_0_RNIKOS1/U0_RGB1_RGB4\ : RGB_NG
      port map(An => \AND2_0_RNIKOS1/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\);
    
    \MemorySynchronizer_0/un1_nreset_31_0_a3\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[3]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_31_i\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[29]\, B => 
        \sb_sb_0_STAMP_PWDATA[29]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[29]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_24\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[24]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_23_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_24_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_24_Z\, 
        CC => NET_CC_CONFIG699, P => NET_CC_CONFIG697, UB => 
        NET_CC_CONFIG698);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_48\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[25]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_48_Z\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_18\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[18]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_17_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_18_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_18_Z\, CC
         => NET_CC_CONFIG779, P => NET_CC_CONFIG777, UB => 
        NET_CC_CONFIG778);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_19\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_20\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_18_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[20]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_19_Z\, CC
         => NET_CC_CONFIG1080, P => NET_CC_CONFIG1078, UB => 
        NET_CC_CONFIG1079);
    
    \STAMP_0/delay_counter_RNIIFLA[12]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \STAMP_0/delay_counter_Z[15]\, B => 
        \STAMP_0/delay_counter_Z[14]\, C => 
        \STAMP_0/delay_counter_Z[13]\, D => 
        \STAMP_0/delay_counter_Z[12]\, Y => 
        \STAMP_0/N_517_i_0_a2_17\);
    
    \MemorySynchronizer_0/un1_nreset_25_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_37\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_25_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_25_rs_Z\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_44_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[28]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_44\);
    
    \STAMP_0/status_async_cycles_2_sqmuxa_0_a3\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/drdy_flank_detected_dms1_0_sqmuxa_1\, 
        B => \STAMP_0/async_state_Z[1]\, C => 
        \STAMP_0/un1_async_prescaler_count\, Y => 
        \STAMP_0/status_async_cycles_2_sqmuxa\);
    
    \MemorySynchronizer_0/resettimercounter[30]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[30]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_6_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[30]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_6\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[6]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[6]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_5\, S => 
        \MemorySynchronizer_0/temp_1[6]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_6\, CC => 
        NET_CC_CONFIG217, P => NET_CC_CONFIG215, UB => 
        NET_CC_CONFIG216);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_84\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[0]\, 
        IPC => OPEN);
    
    \STAMP_0/un45_async_state_cry_5\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \STAMP_0/config_Z[29]\, B => 
        \STAMP_0_data_frame[8]\, C => ADLIB_GND0, D => ADLIB_GND0, 
        FCI => \STAMP_0/un45_async_state_cry_4_Z\, S => OPEN, Y
         => OPEN, FCO => \STAMP_0/un45_async_state_cry_5_FCNET1\, 
        CC => NET_CC_CONFIG531, P => NET_CC_CONFIG529, UB => 
        NET_CC_CONFIG530);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[13]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[13]\, B => 
        \sb_sb_0_Memory_PRDATA[13]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[0]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[0]\, B => 
        \sb_sb_0_Memory_PRDATA[0]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0]\);
    
    \MemorySynchronizer_0/un1_nreset_28_rs_RNIB0RM\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_2538_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[26]\, C => 
        \MemorySynchronizer_0/un1_nreset_28_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[26]\);
    
    \STAMP_0/spi/rx_data[1]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB0_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[1]\);
    
    \MemorySynchronizer_0/TimeStampReg[1]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[1]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[1]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[10]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => \MemorySynchronizer_0/N_1182\, B => 
        \MemorySynchronizer_0/N_2575\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[10]\, D => 
        \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[10]\);
    
    \STAMP_0/PRDATA[23]\ : SLE
      port map(D => \STAMP_0/N_673\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_71\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[23]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_111\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter[0]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[0]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_34_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[0]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg_RNIK90D[21]\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[21]\, B => 
        NN_1, Y => \MemorySynchronizer_0/N_1980_i\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_25_RNIO3CM8\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[27]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[26]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[27]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[26]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[12]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[13]\, CC
         => NET_CC_CONFIG1156, P => NET_CC_CONFIG1154, UB => 
        NET_CC_CONFIG1155);
    
    \MemorySynchronizer_0/SynchStatusReg2[1]\ : SLE
      port map(D => \MemorySynchronizer_0/temp_1[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[1]\);
    
    \MemorySynchronizer_0/un94_in_enable_23\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[15]\, B => 
        \MemorySynchronizer_0/resettimercounter_Z[14]\, C => 
        \MemorySynchronizer_0/resettimercounter_Z[13]\, D => 
        \MemorySynchronizer_0/resettimercounter_Z[0]\, Y => 
        \MemorySynchronizer_0/un94_in_enable_23_Z\);
    
    \STAMP_0/spi/rx_buffer[5]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[5]\);
    
    \STAMP_0/un1_new_avail_0_sqmuxa_2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/un1_new_avail_0_sqmuxa_1\, B => 
        \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_1\, Y => 
        \STAMP_0/un1_new_avail_0_sqmuxa_2_Z\);
    
    \STAMP_0/delay_counter_cry[13]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[13]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[12]\, S
         => \STAMP_0/delay_counter_s[13]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[13]\, CC => NET_CC_CONFIG434, 
        P => NET_CC_CONFIG432, UB => NET_CC_CONFIG433);
    
    \AND2_0_RNIKOS1/U0_RGB1_RGB2\ : RGB_NG
      port map(An => \AND2_0_RNIKOS1/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, YR => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_138\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/numberofnewavails[2]\ : SLE
      port map(D => \MemorySynchronizer_0/ConfigReg_Z[2]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/numberofnewavails_0_sqmuxa\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/numberofnewavails_Z[2]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_180\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA[9]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[9]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[9]\);
    
    \STAMP_0/spi/tx_buffer_RNO[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[1]\, B => 
        \STAMP_0/spi/tx_buffer_Z[0]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_140\);
    
    \MemorySynchronizer_0/N_2538_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_72\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_2538_set_Z\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_35_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_73\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_35_set_Z\);
    
    \STAMP_0/measurement_dms2[6]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[38]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4[13]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \MemorySynchronizer_0/un104_in_enable_13\, B
         => \MemorySynchronizer_0/SynchStatusReg2_Z[13]\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2594\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[13]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_21\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[26]\, B
         => ADLIB_GND0, C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0]\, 
        IPC => OPEN);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.un151_in_enablelto30_15\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/temp_1[13]\, B => 
        \MemorySynchronizer_0/temp_1[14]\, C => 
        \MemorySynchronizer_0/temp_1[15]\, D => 
        \MemorySynchronizer_0/temp_1[16]\, Y => 
        \MemorySynchronizer_0/un151_in_enablelto30_15\);
    
    \MemorySynchronizer_0/un1_nreset_50_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_57_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_50_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_50_rs_Z\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_42_set_RNI0MPP\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_42_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[18]\, C => 
        \MemorySynchronizer_0/un1_nreset_15_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[18]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[5]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_5_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_52\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[21]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[21]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[21]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[21]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[7]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[7]\, 
        B => \sb_sb_0_STAMP_PWDATA[7]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[7]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_0_CC_0\ : 
        CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => CI_TO_CO195, P(0) => 
        ADLIB_VCC1, P(1) => ADLIB_GND0, P(2) => NET_CC_CONFIG197, 
        P(3) => NET_CC_CONFIG200, P(4) => NET_CC_CONFIG203, P(5)
         => NET_CC_CONFIG206, P(6) => NET_CC_CONFIG209, P(7) => 
        NET_CC_CONFIG212, P(8) => NET_CC_CONFIG215, P(9) => 
        NET_CC_CONFIG218, P(10) => NET_CC_CONFIG221, P(11) => 
        NET_CC_CONFIG224, UB(0) => ADLIB_VCC1, UB(1) => 
        ADLIB_GND0, UB(2) => NET_CC_CONFIG198, UB(3) => 
        NET_CC_CONFIG201, UB(4) => NET_CC_CONFIG204, UB(5) => 
        NET_CC_CONFIG207, UB(6) => NET_CC_CONFIG210, UB(7) => 
        NET_CC_CONFIG213, UB(8) => NET_CC_CONFIG216, UB(9) => 
        NET_CC_CONFIG219, UB(10) => NET_CC_CONFIG222, UB(11) => 
        NET_CC_CONFIG225, CC(0) => nc390, CC(1) => nc34, CC(2)
         => NET_CC_CONFIG199, CC(3) => NET_CC_CONFIG202, CC(4)
         => NET_CC_CONFIG205, CC(5) => NET_CC_CONFIG208, CC(6)
         => NET_CC_CONFIG211, CC(7) => NET_CC_CONFIG214, CC(8)
         => NET_CC_CONFIG217, CC(9) => NET_CC_CONFIG220, CC(10)
         => NET_CC_CONFIG223, CC(11) => NET_CC_CONFIG226);
    
    \MemorySynchronizer_0/resettimercounter[4]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[4]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_30_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[4]\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO_0[29]\ : CFG4
      generic map(INIT => x"1030")

      port map(A => \MemorySynchronizer_0/N_2586\, B => 
        \MemorySynchronizer_0/N_2517\, C => 
        \MemorySynchronizer_0/APBState_Z[1]\, D => 
        \sb_sb_0_STAMP_PADDR[4]\, Y => 
        \MemorySynchronizer_0/N_122_i\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[15]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_15\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_0_Z[15]\, 
        C => \MemorySynchronizer_0/N_1213\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[15]\);
    
    \STAMP_0/spi_tx_data_RNO[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[1]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_297_i\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[19]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[19]\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/N_2323\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[19]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[19]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_0\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[0]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => ADLIB_GND0, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_0_Z\, CC
         => NET_CC_CONFIG725, P => NET_CC_CONFIG723, UB => 
        NET_CC_CONFIG724);
    
    \STAMP_0/config[12]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[12]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S[28]\ : 
        CFG4
      generic map(INIT => x"7FFF")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_Z[28]\, B
         => \MemorySynchronizer_0/APBState_Z[0]\, C => 
        \MemorySynchronizer_0/N_271\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_18_0_Z[19]\, Y
         => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[20]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[4]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[20]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[20]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[8]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_60\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[8]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[8]\, D
         => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[8]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[8]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[8]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[25]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[4]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[25]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[25]\);
    
    AFLSDF_INV_20 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_49\, Y => 
        \AFLSDF_INV_20\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_21\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[21]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_20_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_21_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_21_Z\, 
        CC => NET_CC_CONFIG690, P => NET_CC_CONFIG688, UB => 
        NET_CC_CONFIG689);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[26]\ : SLE
      port map(D => \STAMP_0_data_frame[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[26]\);
    
    \LED_HEARTBEAT_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => LED_HEARTBEAT_c, E => ADLIB_VCC1, DOUT => 
        \LED_HEARTBEAT_obuf/U0/DOUT1\, EOUT => 
        \LED_HEARTBEAT_obuf/U0/EOUT1\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_0_CC_1\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO1019, CO => CI_TO_CO1020, P(0) => 
        NET_CC_CONFIG1048, P(1) => NET_CC_CONFIG1051, P(2) => 
        NET_CC_CONFIG1054, P(3) => NET_CC_CONFIG1057, P(4) => 
        NET_CC_CONFIG1060, P(5) => NET_CC_CONFIG1063, P(6) => 
        NET_CC_CONFIG1066, P(7) => NET_CC_CONFIG1069, P(8) => 
        NET_CC_CONFIG1072, P(9) => NET_CC_CONFIG1075, P(10) => 
        NET_CC_CONFIG1078, P(11) => NET_CC_CONFIG1081, UB(0) => 
        NET_CC_CONFIG1049, UB(1) => NET_CC_CONFIG1052, UB(2) => 
        NET_CC_CONFIG1055, UB(3) => NET_CC_CONFIG1058, UB(4) => 
        NET_CC_CONFIG1061, UB(5) => NET_CC_CONFIG1064, UB(6) => 
        NET_CC_CONFIG1067, UB(7) => NET_CC_CONFIG1070, UB(8) => 
        NET_CC_CONFIG1073, UB(9) => NET_CC_CONFIG1076, UB(10) => 
        NET_CC_CONFIG1079, UB(11) => NET_CC_CONFIG1082, CC(0) => 
        NET_CC_CONFIG1050, CC(1) => NET_CC_CONFIG1053, CC(2) => 
        NET_CC_CONFIG1056, CC(3) => NET_CC_CONFIG1059, CC(4) => 
        NET_CC_CONFIG1062, CC(5) => NET_CC_CONFIG1065, CC(6) => 
        NET_CC_CONFIG1068, CC(7) => NET_CC_CONFIG1071, CC(8) => 
        NET_CC_CONFIG1074, CC(9) => NET_CC_CONFIG1077, CC(10) => 
        NET_CC_CONFIG1080, CC(11) => NET_CC_CONFIG1083);
    
    AFLSDF_INV_80 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_80\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[13]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_13\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[27]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[27]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1064\, Y => 
        \MemorySynchronizer_0/N_1095\);
    
    \STAMP_0/spi/sclk_buffer_0_sqmuxa_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/N_30\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/ss_n_buffer_Z[0]\, Y => 
        \STAMP_0/spi/sclk_buffer_0_sqmuxa\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_21\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[23]\, B => 
        \MemorySynchronizer_0/un104_in_enable_22\, C => 
        \MemorySynchronizer_0/un104_in_enable_23\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[22]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[10]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[11]\, CC
         => NET_CC_CONFIG571, P => NET_CC_CONFIG569, UB => 
        NET_CC_CONFIG570);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[18]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_18\);
    
    \MemorySynchronizer_0/un1_nreset_53_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_53\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_53_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_53_rs_Z\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[20]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_20\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[24]\ : SLE
      port map(D => \STAMP_0_data_frame[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[24]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[27]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[27]\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2564\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1411\);
    
    \STAMP_0/measurement_dms1[14]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[62]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[18]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[18]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_29\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un104_in_enable_29\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[29]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_28_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_29_Z\, CC => 
        NET_CC_CONFIG910, P => NET_CC_CONFIG908, UB => 
        NET_CC_CONFIG909);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[11]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_11_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_68\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_103\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[3]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net\, 
        IPC => OPEN);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_13\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/NGMUX1_ARST_N_net\, IPB
         => OPEN, IPC => \sb_sb_0/CCC_0/CCC_INST/PADDR_net[3]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[7]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[7]\, B => 
        \sb_sb_0_STAMP_PWDATA[7]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[7]\);
    
    \STAMP_0/dummy_1_sqmuxa_2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => sb_sb_0_STAMP_PWRITE, B => 
        \STAMP_0/component_state_Z[3]\, C => 
        \sb_sb_0_STAMP_PADDR[9]\, D => \sb_sb_0_STAMP_PADDR[4]\, 
        Y => \STAMP_0/dummy_1_sqmuxa_2_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter[21]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[21]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_43_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[21]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_219\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA[24]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[24]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[24]\);
    
    \STAMP_0/measurement_dms1[11]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[59]\);
    
    AFLSDF_INV_93 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_36_Z\, Y => 
        \AFLSDF_INV_93\);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_19\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[31]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[24]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[23]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[18]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_19_Z\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[5]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_5_S\, 
        Y => \MemorySynchronizer_0/N_1553\);
    
    \MemorySynchronizer_0/un1_nreset_46_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_35\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_46_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_46_rs_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_238\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48]\, 
        IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data_1[18]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[50]\, B => 
        \STAMP_0/dummy_Z[18]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_635\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_15_RNI58K18\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[17]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[16]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[17]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[16]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[7]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[8]\, CC
         => NET_CC_CONFIG1141, P => NET_CC_CONFIG1139, UB => 
        NET_CC_CONFIG1140);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[15]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_15\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_276\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_20\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[20]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_19_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_20_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_20_Z\, 
        CC => NET_CC_CONFIG687, P => NET_CC_CONFIG685, UB => 
        NET_CC_CONFIG686);
    
    \STAMP_0/async_prescaler_count[8]\ : SLE
      port map(D => \STAMP_0/async_prescaler_count_5_Z[8]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[8]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[2]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[2]\, B => 
        \sb_sb_0_Memory_PRDATA[2]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[21]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_21_S\, 
        Y => \MemorySynchronizer_0/N_1497\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_0[3]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[3]\, B => 
        \sb_sb_0_STAMP_PWDATA[3]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_0_Z[3]\);
    
    \STAMP_0/spi/count[3]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[3]\);
    
    \STAMP_0/dummy[19]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_74\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[19]\);
    
    
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_RNIKHI89_FCINST1\ : 
        FCEND_BUFF_CC
      port map(FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_29_RNIKHI89_FCNET1\, 
        CO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[15]\, CC
         => NET_CC_CONFIG1165, P => NET_CC_CONFIG1163, UB => 
        NET_CC_CONFIG1164);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[20]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_20\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[20]\, 
        C => \MemorySynchronizer_0/N_1513\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[20]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_18\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[18]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[18]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_17_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_18_Z\, CC => 
        NET_CC_CONFIG877, P => NET_CC_CONFIG875, UB => 
        NET_CC_CONFIG876);
    
    \STAMP_0/spi/count_lm_0[13]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[13]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[13]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_8\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[8]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[8]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_7_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_8_Z\, CC => 
        NET_CC_CONFIG847, P => NET_CC_CONFIG845, UB => 
        NET_CC_CONFIG846);
    
    \MemorySynchronizer_0/TimeStampGen/un1_prescaler_ac0_5\ : 
        CFG3
      generic map(INIT => x"80")

      port map(A => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[2]\, B => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_c2\, C
         => \MemorySynchronizer_0/TimeStampGen/prescaler_Z[3]\, Y
         => \MemorySynchronizer_0/TimeStampGen/un1_prescaler_c4\);
    
    AFLSDF_INV_96 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_33\, Y => 
        \AFLSDF_INV_96\);
    
    \STAMP_0/config_143_0_0_a3\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \STAMP_0/component_state_Z[5]\, B => 
        \STAMP_0/component_state_Z[3]\, C => \STAMP_0/un76_paddr\, 
        D => sb_sb_0_STAMP_PWRITE, Y => \STAMP_0/config_143\);
    
    \STAMP_0/spi/count_cry[15]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[14]\, S => 
        \STAMP_0/spi/count_s[15]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[15]\, CC => NET_CC_CONFIG970, P
         => NET_CC_CONFIG968, UB => NET_CC_CONFIG969);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[8]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[8]\);
    
    \STAMP_0/async_prescaler_count[10]\ : SLE
      port map(D => \STAMP_0/un5_async_prescaler_count_cry_10_S\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \STAMP_0/async_prescaler_count_Z[10]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[13]\ : SLE
      port map(D => \STAMP_0_data_frame[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[13]\);
    
    \stamp0_spi_clock_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => stamp0_spi_clock_c, E => ADLIB_VCC1, DOUT => 
        \stamp0_spi_clock_obuf/U0/DOUT1\, EOUT => 
        \stamp0_spi_clock_obuf/U0/EOUT1\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[18]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[18]\, B => 
        \sb_sb_0_STAMP_PWDATA[18]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[18]\);
    
    \STAMP_0/un1_spi_rx_data_1[3]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[35]\, B => 
        \STAMP_0/dummy_Z[3]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_620\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_o2_0[19]\ : CFG4
      generic map(INIT => x"0FF8")

      port map(A => \sb_sb_0_STAMP_PADDR[2]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, C => \sb_sb_0_STAMP_PADDR[4]\, 
        D => \sb_sb_0_STAMP_PADDR[5]\, Y => 
        \MemorySynchronizer_0/N_2316\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_272\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_RNIC38O1[0]_CC_0\ : 
        CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => CI_TO_CO1114, P(0) => 
        ADLIB_VCC1, P(1) => ADLIB_VCC1, P(2) => ADLIB_GND0, P(3)
         => NET_CC_CONFIG1115, P(4) => NET_CC_CONFIG1118, P(5)
         => NET_CC_CONFIG1121, P(6) => NET_CC_CONFIG1124, P(7)
         => NET_CC_CONFIG1127, P(8) => NET_CC_CONFIG1130, P(9)
         => NET_CC_CONFIG1133, P(10) => NET_CC_CONFIG1136, P(11)
         => NET_CC_CONFIG1139, UB(0) => ADLIB_VCC1, UB(1) => 
        ADLIB_VCC1, UB(2) => ADLIB_VCC1, UB(3) => 
        NET_CC_CONFIG1116, UB(4) => NET_CC_CONFIG1119, UB(5) => 
        NET_CC_CONFIG1122, UB(6) => NET_CC_CONFIG1125, UB(7) => 
        NET_CC_CONFIG1128, UB(8) => NET_CC_CONFIG1131, UB(9) => 
        NET_CC_CONFIG1134, UB(10) => NET_CC_CONFIG1137, UB(11)
         => NET_CC_CONFIG1140, CC(0) => nc28, CC(1) => nc361, 
        CC(2) => nc115, CC(3) => NET_CC_CONFIG1117, CC(4) => 
        NET_CC_CONFIG1120, CC(5) => NET_CC_CONFIG1123, CC(6) => 
        NET_CC_CONFIG1126, CC(7) => NET_CC_CONFIG1129, CC(8) => 
        NET_CC_CONFIG1132, CC(9) => NET_CC_CONFIG1135, CC(10) => 
        NET_CC_CONFIG1138, CC(11) => NET_CC_CONFIG1141);
    
    \MemorySynchronizer_0/un1_nreset_18_0_a3\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[15]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_18_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_90\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[6]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[18]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[18]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[18]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[18]\);
    
    \STAMP_0/PRDATA[12]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[12]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[13]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[13]\);
    
    \STAMP_0/spi_tx_data_RNO[13]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[13]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_266_i\);
    
    \MemorySynchronizer_0/resynctimercounter[13]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1109\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[13]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL[28]\ : 
        CFG2
      generic map(INIT => x"7")

      port map(A => \MemorySynchronizer_0/N_2595\, B => 
        \MemorySynchronizer_0/APBState_Z[0]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_7\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[7]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_6_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_7_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_7_Z\, CC
         => NET_CC_CONFIG746, P => NET_CC_CONFIG744, UB => 
        NET_CC_CONFIG745);
    
    \STAMP_0/status_async_cycles_lm_0[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/status_async_cycles_3_sqmuxa\, B => 
        \STAMP_0/status_async_cycles_s[2]\, C => 
        \STAMP_0/status_async_cycles_1_sqmuxa_Z\, Y => 
        \STAMP_0/status_async_cycles_lm[2]\);
    
    \STAMP_0/drdy_flank_detected_dms1_0_sqmuxa_1_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \STAMP_0/spi_request_for_Z[1]\, B => 
        \STAMP_0/spi_request_for_Z[0]\, C => 
        \STAMP_0/component_state_Z[0]\, D => \STAMP_0/N_331\, Y
         => \STAMP_0/drdy_flank_detected_dms1_0_sqmuxa_1\);
    
    \STAMP_0/status_async_cycles[0]\ : SLE
      port map(D => \STAMP_0/status_async_cycles_lm[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/status_async_cycles_1_sqmuxa_1_i_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[3]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14[4]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[4]\, 
        B => \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2567\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1265\);
    
    \STAMP_0/spi/count_lm_0[8]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[8]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[8]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[2]\ : SLE
      port map(D => \STAMP_0_data_frame[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[2]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_41\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/ResetTimerValueReg[15]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[15]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[4]\, B => 
        \sb_sb_0_Memory_PRDATA[4]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_19_RNIMMT98\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[21]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[20]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[21]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[20]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[9]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[10]\, CC
         => NET_CC_CONFIG1147, P => NET_CC_CONFIG1145, UB => 
        NET_CC_CONFIG1146);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[10]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[10]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_s_387_CC_2\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO3, CO => OPEN, P(0) => 
        NET_CC_CONFIG67, P(1) => NET_CC_CONFIG70, P(2) => 
        NET_CC_CONFIG73, P(3) => NET_CC_CONFIG76, P(4) => 
        NET_CC_CONFIG79, P(5) => NET_CC_CONFIG82, P(6) => 
        NET_CC_CONFIG85, P(7) => NET_CC_CONFIG88, P(8) => 
        NET_CC_CONFIG91, P(9) => NET_CC_CONFIG94, P(10) => 
        NET_CC_CONFIG97, P(11) => ADLIB_VCC1, UB(0) => 
        NET_CC_CONFIG68, UB(1) => NET_CC_CONFIG71, UB(2) => 
        NET_CC_CONFIG74, UB(3) => NET_CC_CONFIG77, UB(4) => 
        NET_CC_CONFIG80, UB(5) => NET_CC_CONFIG83, UB(6) => 
        NET_CC_CONFIG86, UB(7) => NET_CC_CONFIG89, UB(8) => 
        NET_CC_CONFIG92, UB(9) => NET_CC_CONFIG95, UB(10) => 
        NET_CC_CONFIG98, UB(11) => ADLIB_VCC1, CC(0) => 
        NET_CC_CONFIG69, CC(1) => NET_CC_CONFIG72, CC(2) => 
        NET_CC_CONFIG75, CC(3) => NET_CC_CONFIG78, CC(4) => 
        NET_CC_CONFIG81, CC(5) => NET_CC_CONFIG84, CC(6) => 
        NET_CC_CONFIG87, CC(7) => NET_CC_CONFIG90, CC(8) => 
        NET_CC_CONFIG93, CC(9) => NET_CC_CONFIG96, CC(10) => 
        NET_CC_CONFIG99, CC(11) => nc264);
    
    \MemorySynchronizer_0/ResetTimerValueReg[4]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[4]\);
    
    \STAMP_0/spi/rx_data[4]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB0_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[4]\);
    
    \STAMP_0/config[13]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[13]\);
    
    \STAMP_0/spi/count_lm_0[24]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[24]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[24]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_0_a2_0_0[25]\ : 
        CFG3
      generic map(INIT => x"DC")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[27]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, C
         => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_0_a2_0_0_Z[25]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_124\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6]\, 
        IPC => OPEN);
    
    \STAMP_0/component_state_RNO[1]\ : CFG4
      generic map(INIT => x"BF3F")

      port map(A => \STAMP_0/N_333\, B => \STAMP_0/N_219\, C => 
        \STAMP_0/N_160\, D => \STAMP_0/N_109_i\, Y => 
        \STAMP_0/N_536_i\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_34_set_RNIEN2S\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_34_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[2]\, C
         => \MemorySynchronizer_0/un1_nreset_45_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[2]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[27]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[27]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_29\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[29]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_28_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[3]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_29_Z\, CC
         => NET_CC_CONFIG384, P => NET_CC_CONFIG382, UB => 
        NET_CC_CONFIG383);
    
    AFLSDF_INV_32 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_56_Z\, Y => 
        \AFLSDF_INV_32\);
    
    \STAMP_0/un1_spi_rx_data_2[26]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_609\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, C => \STAMP_0/N_643\, Y
         => \STAMP_0/N_676\);
    
    AFLSDF_INV_101 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_52\, Y => 
        \AFLSDF_INV_101\);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_30\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_25_Z\, 
        B => ENABLE_MEMORY_LED_c, C => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_17_Z\, 
        D => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_16_Z\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_30_Z\);
    
    AFLSDF_INV_2 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_2\);
    
    \MemorySynchronizer_0/waitingtimercounter[16]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[16]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_47_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[16]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[11]\ : SLE
      port map(D => \STAMP_0_data_frame[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[11]\);
    
    AFLSDF_INV_8 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_8\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[24]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[24]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[26]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[24]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_246\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6]\, IPC
         => OPEN);
    
    \MemorySynchronizer_0/un94_in_enable_19\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[30]\, B => 
        \MemorySynchronizer_0/resettimercounter_Z[29]\, C => 
        \MemorySynchronizer_0/resettimercounter_Z[28]\, D => 
        \MemorySynchronizer_0/resettimercounter_Z[27]\, Y => 
        \MemorySynchronizer_0/un94_in_enable_19_Z\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[12]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[12]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1079\, Y => 
        \MemorySynchronizer_0/N_1110\);
    
    \MemorySynchronizer_0/resettimercounter[29]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[29]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_8_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[29]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_11\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[11]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[11]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_10\, S => 
        \MemorySynchronizer_0/temp_1[11]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_11\, CC => 
        NET_CC_CONFIG232, P => NET_CC_CONFIG230, UB => 
        NET_CC_CONFIG231);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[28]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_28_S\, 
        Y => \MemorySynchronizer_0/N_1474\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_57\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[2]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[2]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[2]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[2]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[21]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[21]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[21]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[21]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[21]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[21]\);
    
    \STAMP_0/spi/count[2]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[2]\);
    
    AFLSDF_INV_60 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_60\);
    
    AFLSDF_INV_0 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_41\, Y => 
        \AFLSDF_INV_0\);
    
    \STAMP_0/un1_async_prescaler_countlto5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \STAMP_0/async_prescaler_count_Z[5]\, B => 
        \STAMP_0/async_prescaler_count_Z[4]\, C => 
        \STAMP_0/async_prescaler_count_Z[3]\, D => 
        \STAMP_0/async_prescaler_count_Z[2]\, Y => 
        \STAMP_0/un1_async_prescaler_countlt8\);
    
    \STAMP_0/spi/mosi_cl_RNO\ : CFG4
      generic map(INIT => x"4440")

      port map(A => \STAMP_0/spi/ss_n_buffer_1_sqmuxa\, B => 
        debug_led_net_0, C => mosi_cl, D => 
        \STAMP_0/spi/mosi_1_1_2\, Y => \STAMP_0/spi/N_25_i\);
    
    \STAMP_0/delay_counter_lm_0[25]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[25]\, Y => 
        \STAMP_0/delay_counter_lm[25]\);
    
    \STAMP_0/un1_spi_rx_data_2[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_589\, B => \STAMP_0/N_623\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_656\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[9]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[9]\);
    
    \stamp0_spi_clock_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \stamp0_spi_clock_obuf/U0/DOUT1\, Y => 
        \stamp0_spi_clock_obuf/U0/DOUT\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_109\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1]\, 
        IPB => OPEN, IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_77\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_105\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RCGF_net[5]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[12]\ : SLE
      port map(D => \STAMP_0_data_frame[44]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[12]\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\);
    
    \nCS1_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \nCS1_obuf/U0/DOUT1\, Y => 
        \nCS1_obuf/U0/DOUT\);
    
    \MemorySynchronizer_0/ReadInterrupt\ : SLE
      port map(D => \MemorySynchronizer_0/N_191_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ReadInterrupt_0_sqmuxa_2_i_0_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => MemorySynchronizer_0_ReadInterrupt);
    
    \STAMP_0/PRDATA[1]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[1]\);
    
    \stamp0_ready_temp_ibuf/U0/U_IOINFF\ : IOINFF_BYPASS
      port map(A => \stamp0_ready_temp_ibuf/U0/YIN1\, Y => 
        \stamp0_ready_temp_ibuf/U0/YIN\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_242\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2]\, IPC
         => OPEN);
    
    \MemorySynchronizer_0/TimeStampGen/un6_enable_3\ : CFG4
      generic map(INIT => x"0040")

      port map(A => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[5]\, B => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[4]\, C => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[3]\, D => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[2]\, Y => 
        \MemorySynchronizer_0/TimeStampGen/un6_enable_3_Z\);
    
    \STAMP_0/measurement_dms2[8]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[40]\);
    
    \STAMP_0/delay_counter_lm_0[17]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[17]\, Y => 
        \STAMP_0/delay_counter_lm[17]\);
    
    \MemorySynchronizer_0/PRDATA[25]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[25]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[25]\);
    
    \STAMP_0/spi/clk_toggles_lm_0[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \STAMP_0/spi/ss_n_buffer_1_sqmuxa\, B => 
        \STAMP_0/spi/clk_toggles_Z[0]\, Y => 
        \STAMP_0/spi/clk_toggles_lm[0]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[3]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[3]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[1]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[1]\, B => 
        \sb_sb_0_STAMP_PWDATA[1]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[1]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[12]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[12]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0[4]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/N_1265\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[4]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[4]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[4]\, Y => 
        \MemorySynchronizer_0/PRDATA_21[4]\);
    
    \MemorySynchronizer_0/un1_nreset_14\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[19]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_14_i\);
    
    \STAMP_0/measurement_dms1[13]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[61]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[14]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[14]\, B => 
        \sb_sb_0_Memory_PRDATA[14]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[27]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_27_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[5]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[9]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[9]\, B => 
        \sb_sb_0_STAMP_PWDATA[9]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[9]\);
    
    \MemorySynchronizer_0/un1_nreset_35_rs_RNIT83G\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_42_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[30]\, C
         => \MemorySynchronizer_0/un1_nreset_35_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[30]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_160\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_154\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_28\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_29\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_27_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[29]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_28_Z\, CC
         => NET_CC_CONFIG1107, P => NET_CC_CONFIG1105, UB => 
        NET_CC_CONFIG1106);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[12]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[12]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[12]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[12]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[24]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[24]\, B => 
        \MemorySynchronizer_0/un104_in_enable_24\, C => 
        \MemorySynchronizer_0/N_2574\, D => 
        \MemorySynchronizer_0/N_2577\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[24]\);
    
    \MemorySynchronizer_0/un1_nreset_16\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[17]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_16_i\);
    
    \STAMP_0/dummy[10]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_75\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[10]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[19]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[19]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4[6]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \MemorySynchronizer_0/un104_in_enable_6\, B
         => \MemorySynchronizer_0/SynchStatusReg2_Z[6]\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2594\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[6]\);
    
    \STAMP_0/async_state_17_iv_0[1]\ : CFG4
      generic map(INIT => x"FF41")

      port map(A => \STAMP_0/un1_async_state_0_sqmuxa_i\, B => 
        \STAMP_0/N_206\, C => \STAMP_0/async_state_Z[1]\, D => 
        \STAMP_0/request_resync_1_sqmuxa_1_Z\, Y => 
        \STAMP_0/async_state_17[1]\);
    
    \STAMP_0/PRDATA[19]\ : SLE
      port map(D => \STAMP_0/N_669\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_76\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[19]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_271\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net\, 
        IPC => OPEN);
    
    \STAMP_0/un1_component_state_14_i_o2_RNO\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => \STAMP_0/drdy_flank_detected_dms1_Z\, B => 
        \STAMP_0/config_Z[30]\, C => 
        \STAMP_0/component_state_Z[5]\, D => \STAMP_0/N_238\, Y
         => \STAMP_0/N_110_i\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[21]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[21]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1070\, Y => 
        \MemorySynchronizer_0/N_1101\);
    
    \STAMP_0/un52_paddr_2_0\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \sb_sb_0_STAMP_PADDR[0]\, B => 
        \sb_sb_0_STAMP_PADDR[1]\, C => \sb_sb_0_STAMP_PADDR[6]\, 
        D => \sb_sb_0_STAMP_PADDR[5]\, Y => 
        \STAMP_0/un52_paddr_2_0_Z\);
    
    \STAMP_0/spi/sclk_buffer\ : SLE
      port map(D => \STAMP_0/spi/N_20_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        debug_led_net_0, ALn => ADLIB_VCC1, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => stamp0_spi_clock_c);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[29]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[29]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[29]\, C => 
        \MemorySynchronizer_0/N_2598\, D => 
        \MemorySynchronizer_0/N_2576\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[29]\);
    
    \MemorySynchronizer_0/TimeStampReg[2]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[2]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampReg_Z[2]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[30]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[30]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[30]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_60\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[7]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[7]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1084\, Y => 
        \MemorySynchronizer_0/N_1115\);
    
    \STAMP_0/component_state_ns_i_0_a2[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \STAMP_0/N_238\, B => \STAMP_0/spi_busy\, Y
         => \STAMP_0/N_331\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_106\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net\, IPC
         => OPEN);
    
    \STAMP_0/spi/rx_data[5]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[5]\);
    
    \STAMP_0/spi/tx_buffer_RNO[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[4]\, B => 
        \STAMP_0/spi/tx_buffer_Z[3]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_134\);
    
    \STAMP_0/spi/rx_buffer[13]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[13]\);
    
    \STAMP_0/spi/count_cry[14]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[14]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[13]\, S => 
        \STAMP_0/spi/count_s[14]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[14]\, CC => NET_CC_CONFIG967, P
         => NET_CC_CONFIG965, UB => NET_CC_CONFIG966);
    
    \MemorySynchronizer_0/waitingtimercounter_RNI2T2L[21]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_39_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[21]\, C
         => \MemorySynchronizer_0/un1_nreset_43_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[21]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_29\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[29]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_28_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_29_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_29_Z\, CC
         => NET_CC_CONFIG812, P => NET_CC_CONFIG810, UB => 
        NET_CC_CONFIG811);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_204\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_GND0, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_RNO[5]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[5]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, C
         => \MemorySynchronizer_0/SynchStatusReg_Z[7]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_m[7]\);
    
    \STAMP_0/spi/count[29]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[29]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB12_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[29]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[22]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_22\);
    
    \MemorySynchronizer_0/PRDATA[28]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[28]\);
    
    \STAMP_0/un1_spi_rx_data_2[14]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_597\, B => \STAMP_0/N_631\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_664\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[20]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[20]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_37\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[23]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_37_Z\);
    
    \MemorySynchronizer_0/MemorySyncState[2]\ : SLE
      port map(D => \MemorySynchronizer_0/N_304\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        ENABLE_MEMORY_LED_c, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/MemorySyncState_Z[2]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_54\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_25\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[25]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_24_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_25_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_25_Z\, 
        CC => NET_CC_CONFIG702, P => NET_CC_CONFIG700, UB => 
        NET_CC_CONFIG701);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[21]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[21]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[20]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[21]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[21]\, CC
         => NET_CC_CONFIG69, P => NET_CC_CONFIG67, UB => 
        NET_CC_CONFIG68);
    
    \MemorySynchronizer_0/PRDATA[1]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[1]\);
    
    \STAMP_0/delay_counter[9]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[9]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_4\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[4]\, 
        B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_3_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_4_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_4_Z\, 
        CC => NET_CC_CONFIG639, P => NET_CC_CONFIG637, UB => 
        NET_CC_CONFIG638);
    
    \MemorySynchronizer_0/un1_nreset_38_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[27]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_38_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_74\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[30]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[30]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_30\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_113\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_28\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[28]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[28]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_27\, S => 
        \MemorySynchronizer_0/temp_1[28]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_28\, CC => 
        NET_CC_CONFIG283, P => NET_CC_CONFIG281, UB => 
        NET_CC_CONFIG282);
    
    \MemorySynchronizer_0/un1_nreset_52_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_52\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_52_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_52_rs_Z\);
    
    \STAMP_0/spi/rx_data[15]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[15]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_12\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[12]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_11_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_12_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_12_Z\, 
        CC => NET_CC_CONFIG663, P => NET_CC_CONFIG661, UB => 
        NET_CC_CONFIG662);
    
    \STAMP_0/measurement_temp[15]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[31]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_89\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[5]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un104_in_enable_cry_24\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un104_in_enable_24\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[24]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_23_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_24_Z\, CC => 
        NET_CC_CONFIG895, P => NET_CC_CONFIG893, UB => 
        NET_CC_CONFIG894);
    
    \STAMP_0/un1_spi_rx_data_2[29]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_612\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, C => \STAMP_0/N_646\, Y
         => \STAMP_0/N_679\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_38_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[15]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_38\);
    
    \STAMP_0/spi/un10_count_0_a2_0_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \STAMP_0/spi/clk_toggles_Z[2]\, B => 
        \STAMP_0/spi/clk_toggles_Z[3]\, Y => 
        \STAMP_0/spi/un10_count_0_a2_0_0_Z\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_5\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[5]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[5]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_4_Z\, S => OPEN, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_5_Z\, CC => 
        NET_CC_CONFIG838, P => NET_CC_CONFIG836, UB => 
        NET_CC_CONFIG837);
    
    \STAMP_0/delay_counter_lm_0[23]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[23]\, Y => 
        \STAMP_0/delay_counter_lm[23]\);
    
    \MemorySynchronizer_0/un1_nreset_28_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_47_i_i_a2_Z\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_28_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_28_rs_Z\);
    
    \STAMP_0/spi_tx_data_RNO[4]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[4]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_294_i\);
    
    \stamp0_spi_dms1_cs_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \stamp0_spi_dms1_cs_obuf/U0/DOUT1\, Y => 
        \stamp0_spi_dms1_cs_obuf/U0/DOUT\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[23]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_23\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[23]\, 
        C => \MemorySynchronizer_0/N_1505\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[23]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[22]\ : SLE
      port map(D => \STAMP_0_data_frame[22]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[22]\);
    
    \STAMP_0/delay_counter_cry[26]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[26]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[25]\, S
         => \STAMP_0/delay_counter_s[26]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[26]\, CC => NET_CC_CONFIG473, 
        P => NET_CC_CONFIG471, UB => NET_CC_CONFIG472);
    
    \STAMP_0/PRDATA[30]\ : SLE
      port map(D => \STAMP_0/N_119_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[30]\);
    
    \MemorySynchronizer_0/waitingtimercounter_RNIR41V[20]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_32_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[20]\, C
         => \MemorySynchronizer_0/un1_nreset_62_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[20]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_32_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_77\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_32_set_Z\);
    
    \STAMP_0/async_state_1_sqmuxa_i_o3\ : CFG4
      generic map(INIT => x"10FF")

      port map(A => \STAMP_0/spi_request_for_Z[1]\, B => 
        \STAMP_0/async_state_Z[1]\, C => \STAMP_0/N_331\, D => 
        \STAMP_0/component_state_Z[0]\, Y => \STAMP_0/N_197\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_28\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[28]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_27_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[4]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_28_Z\, CC
         => NET_CC_CONFIG381, P => NET_CC_CONFIG379, UB => 
        NET_CC_CONFIG380);
    
    \STAMP_0/delay_counter_cry[14]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[14]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[13]\, S
         => \STAMP_0/delay_counter_s[14]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[14]\, CC => NET_CC_CONFIG437, 
        P => NET_CC_CONFIG435, UB => NET_CC_CONFIG436);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_61_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[17]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_61\);
    
    \STAMP_0/spi_dms2_cs_13_iv_i\ : CFG3
      generic map(INIT => x"13")

      port map(A => \STAMP_0/component_state_Z[3]\, B => 
        \STAMP_0/spi_dms2_cs_1_sqmuxa_1\, C => 
        \sb_sb_0_STAMP_PADDR[5]\, Y => 
        \STAMP_0/spi_dms2_cs_13_iv_i_Z\);
    
    AFLSDF_INV_6 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_53_i_i_a2_Z\, 
        Y => \AFLSDF_INV_6\);
    
    \sb_sb_0/Memory_0_intr_or_0\ : CFG3
      generic map(INIT => x"fe")

      port map(A => MemorySynchronizer_0_SynchronizerInterrupt, B
         => MemorySynchronizer_0_ReadInterrupt, C => ADLIB_GND0, 
        Y => \sb_sb_0/Memory_0_intr_or_0_Y\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[26]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[26]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[26]\, D
         => \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[26]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_9[5]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \MemorySynchronizer_0/N_2567\, B => 
        \MemorySynchronizer_0/N_271\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[5]\, D => 
        \sb_sb_0_STAMP_PADDR[6]\, Y => 
        \MemorySynchronizer_0/N_1365\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[14]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[14]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[14]\, C => 
        \MemorySynchronizer_0/N_2598\, D => 
        \MemorySynchronizer_0/N_2576\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[14]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[29]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_29_S\, 
        Y => \MemorySynchronizer_0/N_1480\);
    
    AND2_0_RNIKOS1 : GB_NG
      port map(An => \AFLSDF_INV_78\, ENn => ADLIB_GND0, YNn => 
        \AND2_0_RNIKOS1/U0_YNn\, YSn => 
        \AND2_0_RNIKOS1/U0_YNn_GSouth\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_59\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[13]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_59_Z\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_0_CC_2\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO294, CO => OPEN, P(0) => 
        NET_CC_CONFIG367, P(1) => NET_CC_CONFIG370, P(2) => 
        NET_CC_CONFIG373, P(3) => NET_CC_CONFIG376, P(4) => 
        NET_CC_CONFIG379, P(5) => NET_CC_CONFIG382, P(6) => 
        NET_CC_CONFIG385, P(7) => NET_CC_CONFIG388, P(8) => 
        ADLIB_VCC1, P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, 
        P(11) => ADLIB_VCC1, UB(0) => NET_CC_CONFIG368, UB(1) => 
        NET_CC_CONFIG371, UB(2) => NET_CC_CONFIG374, UB(3) => 
        NET_CC_CONFIG377, UB(4) => NET_CC_CONFIG380, UB(5) => 
        NET_CC_CONFIG383, UB(6) => NET_CC_CONFIG386, UB(7) => 
        NET_CC_CONFIG389, UB(8) => ADLIB_VCC1, UB(9) => 
        ADLIB_VCC1, UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, 
        CC(0) => NET_CC_CONFIG369, CC(1) => NET_CC_CONFIG372, 
        CC(2) => NET_CC_CONFIG375, CC(3) => NET_CC_CONFIG378, 
        CC(4) => NET_CC_CONFIG381, CC(5) => NET_CC_CONFIG384, 
        CC(6) => NET_CC_CONFIG387, CC(7) => NET_CC_CONFIG390, 
        CC(8) => nc398, CC(9) => nc192, CC(10) => nc319, CC(11)
         => nc134);
    
    \STAMP_0/spi/count[17]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[17]\);
    
    \MemorySynchronizer_0/end_one_counter[0]\ : SLE
      port map(D => \MemorySynchronizer_0/N_207_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => ADLIB_VCC1, ADn => ADLIB_VCC1, SLn => 
        ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/end_one_counter_Z[0]\);
    
    \adc_start_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => adc_start_c, E => ADLIB_VCC1, DOUT => 
        \adc_start_obuf/U0/DOUT1\, EOUT => 
        \adc_start_obuf/U0/EOUT1\);
    
    \STAMP_0/un5_async_prescaler_count_cry_8\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[8]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_7_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_8_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_8_Z\, CC
         => NET_CC_CONFIG504, P => NET_CC_CONFIG502, UB => 
        NET_CC_CONFIG503);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_20\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[29]\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[25]\, C => 
        \MemorySynchronizer_0/waitingtimercounter_Z[24]\, D => 
        \MemorySynchronizer_0/waitingtimercounter_Z[22]\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_20_Z\);
    
    \STAMP_0/spi/count_lm_0[12]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[12]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[12]\);
    
    \STAMP_0/measurement_dms1[5]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[53]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_241\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_GND0, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1]\, IPC
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_BREADY_net\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_RNO[19]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_19_S\, 
        Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[12]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[17]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[17]\, B => 
        \sb_sb_0_STAMP_PWDATA[17]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[17]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[30]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[30]\, C => 
        \MemorySynchronizer_0/N_2596\, D => 
        \MemorySynchronizer_0/N_2595\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[30]\);
    
    AFLSDF_INV_79 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_59\, Y => 
        \AFLSDF_INV_79\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_33\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[8]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_ResetTimerValueReg_33_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[0]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[0]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[2]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[0]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_32_i_i_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[28]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_32_i_i_a2_Z\);
    
    \STAMP_0/component_state_ns_0_a3_2_a2[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => sb_sb_0_STAMP_PENABLE, B => 
        \STAMP_0/component_state_Z[4]\, Y => 
        \STAMP_0/apb_spi_finished_0_sqmuxa\);
    
    \STAMP_0/un1_spi_rx_data_0[16]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[16]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[16]\, Y
         => \STAMP_0/N_599\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_91\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[7]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_43_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[21]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_43_i\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_6\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[6]\, 
        B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_5_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_6_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_6_Z\, 
        CC => NET_CC_CONFIG645, P => NET_CC_CONFIG643, UB => 
        NET_CC_CONFIG644);
    
    \MemorySynchronizer_0/ResetTimerValueReg[31]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[31]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[31]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[29]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[29]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[29]\);
    
    AFLSDF_INV_77 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_32\, Y => 
        \AFLSDF_INV_77\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_11\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[11]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_10_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_11_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_11_Z\, CC
         => NET_CC_CONFIG758, P => NET_CC_CONFIG756, UB => 
        NET_CC_CONFIG757);
    
    \STAMP_0/spi/rx_data[11]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[11]\);
    
    \MemorySynchronizer_0/resettimercounter[8]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[8]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_61_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[8]\);
    
    \MemorySynchronizer_0/un1_nreset_5_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_36\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_5_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_5_rs_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO[31]\ : CFG4
      generic map(INIT => x"00AE")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[31]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_152_ss0_i_0\, C
         => \MemorySynchronizer_0/SynchStatusReg_152_sm0\, D => 
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa\, Y
         => \MemorySynchronizer_0/N_2016_i\);
    
    \STAMP_0/un1_spi_rx_data_2[27]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_610\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, C => \STAMP_0/N_644\, Y
         => \STAMP_0/N_677\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_12\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[12]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[12]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_11\, S => 
        \MemorySynchronizer_0/temp_1[12]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_12\, CC => 
        NET_CC_CONFIG235, P => NET_CC_CONFIG233, UB => 
        NET_CC_CONFIG234);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[8]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_8_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_60\);
    
    \STAMP_0/delay_counter[7]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[7]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[21]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[21]\);
    
    \MemorySynchronizer_0/PRDATA[21]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[21]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[21]\);
    
    \STAMP_0/config[27]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[27]\);
    
    \STAMP_0/un1_spi_rx_data[15]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_665\, C => \STAMP_0/spi_rx_data[15]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[15]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_59_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_79\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_59_set_Z\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_38_set_RNISO8K\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_38_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[22]\, C => 
        \MemorySynchronizer_0/un1_nreset_11_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[22]\);
    
    \STAMP_0/PRDATA[22]\ : SLE
      port map(D => \STAMP_0/N_672\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_80\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[22]\);
    
    \MemorySynchronizer_0/resettimercounter[15]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_18_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[15]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_200\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg2_RNO[23]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[2]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[23]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[23]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_16[19]\ : CFG3
      generic map(INIT => x"80")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_18_0_Z[19]\, B
         => \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[2]\, Y => 
        \MemorySynchronizer_0/N_2598\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_22[10]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \sb_sb_0_STAMP_PADDR[5]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, C => 
        \MemorySynchronizer_0/N_271\, D => 
        \MemorySynchronizer_0/N_2564\, Y => 
        \MemorySynchronizer_0/N_2576\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[0]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_0\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[0]\, 
        C => \MemorySynchronizer_0/N_1557\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[0]\);
    
    \STAMP_0/spi/count[6]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[6]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_20\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[20]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[20]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_19_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_20_Z\, CC => 
        NET_CC_CONFIG883, P => NET_CC_CONFIG881, UB => 
        NET_CC_CONFIG882);
    
    \STAMP_0/delay_counter_cry[22]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[22]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[21]\, S
         => \STAMP_0/delay_counter_s[22]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[22]\, CC => NET_CC_CONFIG461, 
        P => NET_CC_CONFIG459, UB => NET_CC_CONFIG460);
    
    \STAMP_0/measurement_dms1[15]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[63]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[8]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => \MemorySynchronizer_0/N_2597\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[8]\, C => 
        \MemorySynchronizer_0/TimeStampReg_Z[8]\, D => 
        \MemorySynchronizer_0/N_1245\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[8]\);
    
    \MemorySynchronizer_0/ConfigReg[28]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[28]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[3]\ : SLE
      port map(D => \STAMP_0_data_frame[35]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[3]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[11]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[11]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[13]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[11]\);
    
    \STAMP_0/spi/count_cry[16]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[16]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[15]\, S => 
        \STAMP_0/spi/count_s[16]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[16]\, CC => NET_CC_CONFIG973, P
         => NET_CC_CONFIG971, UB => NET_CC_CONFIG972);
    
    \MemorySynchronizer_0/un1_nreset_59_rs_RNIVA8U\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_59_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[7]\, C
         => \MemorySynchronizer_0/un1_nreset_59_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[7]\);
    
    \STAMP_0/un5_async_prescaler_count_cry_1\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[1]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_s_1_391_FCO\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_1_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_1_Z\, CC
         => NET_CC_CONFIG483, P => NET_CC_CONFIG481, UB => 
        NET_CC_CONFIG482);
    
    \MemorySynchronizer_0/TimeStampGen/counter[30]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[30]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[30]\);
    
    \MemorySynchronizer_0/TimeStampReg[28]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[28]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[28]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[24]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[24]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[2]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[2]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[2]\, D => 
        \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[2]\);
    
    \MemorySynchronizer_0/numberofnewavails_RNIEAMF1[0]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[2]\, 
        B => \MemorySynchronizer_0/numberofnewavails_Z[1]\, C => 
        \MemorySynchronizer_0/numberofnewavails_Z[0]\, D => 
        \MemorySynchronizer_0/N_140_1_i\, Y => 
        \MemorySynchronizer_0/numberofnewavails_RNIEAMF1_Z[0]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_1_0[10]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[10]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[10]\, C => 
        \MemorySynchronizer_0/N_2576\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[10]\);
    
    \MemorySynchronizer_0/resynctimercounter[21]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1101\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[21]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[11]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_11\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[11]\, 
        C => \MemorySynchronizer_0/N_1537\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[11]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[25]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_25_S\, 
        Y => \MemorySynchronizer_0/N_2422\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_57\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[5]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_ResetTimerValueReg_57_Z\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[11]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[11]\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_9\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/PLL_BYPASS_N_net\, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX3_SEL_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[7]\);
    
    \STAMP_0/PRDATA[5]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[5]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[18]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[2]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[18]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[18]\);
    
    \MemorySynchronizer_0/waitingtimercounter[31]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[31]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_axb_31\);
    
    \MemorySynchronizer_0/un1_nreset_51_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[15]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_51_i\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_18\ : CFG4
      generic map(INIT => x"0002")

      port map(A => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_1_Z\, B
         => \MemorySynchronizer_0/N_1091\, C => 
        \MemorySynchronizer_0/N_1080\, D => 
        \MemorySynchronizer_0/N_1064\, Y => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_18_Z\);
    
    \STAMP_0/spi_tx_data[7]\ : SLE
      port map(D => \STAMP_0/N_291_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[7]\);
    
    \STAMP_0/drdy_flank_detected_dms2_RNIK45E1\ : CFG4
      generic map(INIT => x"FE00")

      port map(A => \STAMP_0/drdy_flank_detected_dms2_Z\, B => 
        \STAMP_0/drdy_flank_detected_temp_Z\, C => 
        \STAMP_0/drdy_flank_detected_dms1_Z\, D => 
        \STAMP_0/config_Z[30]\, Y => \STAMP_0/N_109_i\);
    
    \stamp0_ready_dms2_ibuf/U0/U_IOIN\ : IOIN_IB
      port map(YIN => \stamp0_ready_dms2_ibuf/U0/YIN\, E => 
        ADLIB_GND0, Y => stamp0_ready_dms2_c);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_119\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net\, IPC
         => OPEN);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[14]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[14]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1077\, Y => 
        \MemorySynchronizer_0/N_1108\);
    
    \MemorySynchronizer_0/numberofpendingresyncrequest[2]\ : SLE
      port map(D => \MemorySynchronizer_0/ConfigReg_Z[6]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => \MemorySynchronizer_0/numberofnewavails_0_sqmuxa\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/numberofpendingresyncrequest_Z[2]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_31\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_axb_31\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_30_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_31_FCNET1\, CC
         => NET_CC_CONFIG916, P => NET_CC_CONFIG914, UB => 
        NET_CC_CONFIG915);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_115\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[1]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_1_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[31]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[13]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, B
         => \MemorySynchronizer_0/resettimercounter_Z[13]\, Y => 
        \MemorySynchronizer_0/resettimercounter_m[13]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_7_1[31]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_2561\, C => 
        \sb_sb_0_STAMP_PADDR[2]\, Y => 
        \MemorySynchronizer_0/N_1204_1\);
    
    \sb_sb_0/SYSRESET_POR/IP_INTERFACE_0\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/SYSRESET_POR/UTDO_net\, IPB => OPEN, IPC
         => OPEN);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_1\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[1]\, 
        B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_1_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_1_Z\, 
        CC => NET_CC_CONFIG630, P => NET_CC_CONFIG628, UB => 
        NET_CC_CONFIG629);
    
    \STAMP_0/spi/un10_count_0_a2_RNI2V9I1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \STAMP_0/spi/un7_count_NE_i\, B => 
        \STAMP_0/spi/state_Z[0]\, C => \STAMP_0/spi/un10_count_i\, 
        Y => \STAMP_0/spi/N_50_i\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0_CC_1\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO623, CO => CI_TO_CO624, P(0) => 
        NET_CC_CONFIG658, P(1) => NET_CC_CONFIG661, P(2) => 
        NET_CC_CONFIG664, P(3) => NET_CC_CONFIG667, P(4) => 
        NET_CC_CONFIG670, P(5) => NET_CC_CONFIG673, P(6) => 
        NET_CC_CONFIG676, P(7) => NET_CC_CONFIG679, P(8) => 
        NET_CC_CONFIG682, P(9) => NET_CC_CONFIG685, P(10) => 
        NET_CC_CONFIG688, P(11) => NET_CC_CONFIG691, UB(0) => 
        NET_CC_CONFIG659, UB(1) => NET_CC_CONFIG662, UB(2) => 
        NET_CC_CONFIG665, UB(3) => NET_CC_CONFIG668, UB(4) => 
        NET_CC_CONFIG671, UB(5) => NET_CC_CONFIG674, UB(6) => 
        NET_CC_CONFIG677, UB(7) => NET_CC_CONFIG680, UB(8) => 
        NET_CC_CONFIG683, UB(9) => NET_CC_CONFIG686, UB(10) => 
        NET_CC_CONFIG689, UB(11) => NET_CC_CONFIG692, CC(0) => 
        NET_CC_CONFIG660, CC(1) => NET_CC_CONFIG663, CC(2) => 
        NET_CC_CONFIG666, CC(3) => NET_CC_CONFIG669, CC(4) => 
        NET_CC_CONFIG672, CC(5) => NET_CC_CONFIG675, CC(6) => 
        NET_CC_CONFIG678, CC(7) => NET_CC_CONFIG681, CC(8) => 
        NET_CC_CONFIG684, CC(9) => NET_CC_CONFIG687, CC(10) => 
        NET_CC_CONFIG690, CC(11) => NET_CC_CONFIG693);
    
    \sb_sb_0/FABOSC_0/I_RCOSC_25_50MHZ\ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.000000)

      port map(CLKOUT => 
        \sb_sb_0/FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC\);
    
    \STAMP_0/spi/un10_count_0_a2_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \STAMP_0/spi/clk_toggles_Z[1]\, B => 
        \STAMP_0/spi/clk_toggles_Z[4]\, Y => 
        \STAMP_0/spi/un10_count_0_a2_0_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[11]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[11]\, B => 
        \MemorySynchronizer_0/un104_in_enable_11\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[11]\);
    
    \STAMP_0/un1_spi_rx_data_1[24]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[56]\, B => 
        \STAMP_0/dummy_Z[24]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_641\);
    
    \MemorySynchronizer_0/ConfigReg[31]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[31]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[31]\);
    
    \STAMP_0/PRDATA[2]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[2]\);
    
    \MemorySynchronizer_0/un1_nreset_21\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[13]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_21_i\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_6\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/CLK2_net\, IPB => OPEN, 
        IPC => \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[4]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[29]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[29]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[28]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[29]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[29]\, CC
         => NET_CC_CONFIG93, P => NET_CC_CONFIG91, UB => 
        NET_CC_CONFIG92);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[29]\, B => 
        \sb_sb_0_Memory_PRDATA[29]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[29]\);
    
    \STAMP_0/component_state_RNIFR114[0]\ : CFG3
      generic map(INIT => x"CD")

      port map(A => \STAMP_0/component_state_Z[5]\, B => 
        \STAMP_0/N_238\, C => \STAMP_0/component_state_Z[0]\, Y
         => \STAMP_0/component_state_RNIFR114_Z[0]\);
    
    \STAMP_0/dummy[29]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[29]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_81\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[29]\);
    
    \MemorySynchronizer_0/TimeStampReg[18]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[18]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[18]\);
    
    \STAMP_0/component_state_ns_0_0[1]\ : CFG4
      generic map(INIT => x"AEAA")

      port map(A => \STAMP_0/component_state_ns_0_0_0_Z[1]\, B
         => sb_sb_0_STAMP_PSELx, C => \STAMP_0/N_109_i\, D => 
        \STAMP_0/N_333\, Y => \STAMP_0/component_state_ns[1]\);
    
    \MemorySynchronizer_0/un94_in_enable_22\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[12]\, B => 
        \MemorySynchronizer_0/resettimercounter_Z[11]\, C => 
        \MemorySynchronizer_0/resettimercounter_Z[10]\, D => 
        \MemorySynchronizer_0/resettimercounter_Z[9]\, Y => 
        \MemorySynchronizer_0/un94_in_enable_22_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[9]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[9]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[9]\, D => 
        \MemorySynchronizer_0/un5_resettimercounter_m[23]\, Y => 
        \MemorySynchronizer_0/resettimercounter_9[9]\);
    
    \MemorySynchronizer_0/N_2534_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_82\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_2534_set_Z\);
    
    \MemorySynchronizer_0/un1_nreset_54_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_54\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_54_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_54_rs_Z\);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[25]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[25]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1066\, Y => 
        \MemorySynchronizer_0/N_1097\);
    
    \MemorySynchronizer_0/resynceventpulldowncounter_RNO[2]\ : 
        CFG4
      generic map(INIT => x"AA6A")

      port map(A => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[2]\, B
         => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[1]\, C
         => 
        \MemorySynchronizer_0/resynceventpulldowncounter_Z[0]\, D
         => \MemorySynchronizer_0/N_2333\, Y => 
        \MemorySynchronizer_0/N_1052_i_i\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[10]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[10]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[10]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[10]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[10]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[10]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[20]\ : SLE
      port map(D => \STAMP_0_data_frame[52]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[20]\);
    
    \STAMP_0/spi_temp_cs\ : SLE
      port map(D => \STAMP_0/spi_temp_cs_13_iv_i_Z\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_component_state_13_i_0_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => stamp0_spi_temp_cs_c);
    
    \STAMP_0/spi/rx_data[9]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[9]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_13\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_14\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_12_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[14]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_13_Z\, CC
         => NET_CC_CONFIG1062, P => NET_CC_CONFIG1060, UB => 
        NET_CC_CONFIG1061);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[25]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_25\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[25]\, 
        C => \MemorySynchronizer_0/N_2422\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[25]\);
    
    \MemorySynchronizer_0/waitingtimercounter[22]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[22]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_22_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[22]\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0_a3_0_a2[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[1]\, 
        B => \MemorySynchronizer_0/end_one_counter_Z[1]\, Y => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa\);
    
    \MemorySynchronizer_0/APBState_ns_1_0_.m5_0_a3_0_a2\ : CFG4
      generic map(INIT => x"0800")

      port map(A => sb_sb_0_STAMP_PENABLE, B => 
        sb_sb_0_Memory_PSELx, C => \MemorySynchronizer_0/N_301\, 
        D => sb_sb_0_STAMP_PWRITE, Y => 
        \MemorySynchronizer_0/APBState_ns[1]\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => OPEN, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_41_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[4]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_41\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_RNO[17]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_17_S\, 
        Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[14]\);
    
    \STAMP_0/spi/count_cry[3]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[3]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[2]\, S => 
        \STAMP_0/spi/count_s[3]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[3]\, CC => NET_CC_CONFIG934, P
         => NET_CC_CONFIG932, UB => NET_CC_CONFIG933);
    
    \STAMP_0/measurement_temp_1_sqmuxa_0_a3\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \STAMP_0/apb_spi_finished_0_sqmuxa_1\, B => 
        debug_led_net_0, C => \STAMP_0/spi_request_for_Z[1]\, D
         => \STAMP_0/spi_request_for_Z[0]\, Y => 
        \STAMP_0/measurement_temp_1_sqmuxa\);
    
    \MemorySynchronizer_0/un1_nreset_36_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[29]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_36_i\);
    
    \STAMP_0/un1_spi_rx_data_0[19]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[19]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[19]\, Y
         => \STAMP_0/N_602\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_61\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un104_in_enable_cry_27\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un104_in_enable_27\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[27]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_26_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_27_Z\, CC => 
        NET_CC_CONFIG904, P => NET_CC_CONFIG902, UB => 
        NET_CC_CONFIG903);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[14]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[14]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[13]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[14]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[14]\, CC
         => NET_CC_CONFIG48, P => NET_CC_CONFIG46, UB => 
        NET_CC_CONFIG47);
    
    \MemorySynchronizer_0/TimeStampGen/prescaler[5]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc5_Z\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[5]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[15]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[15]\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/N_2323\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[15]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[15]\);
    
    \MemorySynchronizer_0/un1_nreset_12_0_a3\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[21]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_12_i\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_13\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[13]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_12_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[19]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_13_Z\, CC
         => NET_CC_CONFIG336, P => NET_CC_CONFIG334, UB => 
        NET_CC_CONFIG335);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_116\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_10_rs_RNIRIVU\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_37_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[23]\, C => 
        \MemorySynchronizer_0/un1_nreset_10_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[23]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_0_a1\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_0_a1_1_Z\, 
        B => \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[5]\, D => 
        \MemorySynchronizer_0/N_2569\, Y => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_0_a1_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[26]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[26]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[26]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[26]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_0\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[0]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[0]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => ADLIB_GND0, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_0_Z\, CC => 
        NET_CC_CONFIG823, P => NET_CC_CONFIG821, UB => 
        NET_CC_CONFIG822);
    
    \STAMP_0/un1_spi_rx_data[13]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_663\, C => \STAMP_0/spi_rx_data[13]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[13]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[18]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[18]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[18]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_58_i_i_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[8]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_58_i_i_a2_Z\);
    
    \STAMP_0/un1_component_state_13_i_a2_1\ : CFG2
      generic map(INIT => x"2")

      port map(A => \STAMP_0/N_337\, B => 
        \STAMP_0/component_state_Z[0]\, Y => \STAMP_0/N_364\);
    
    \STAMP_0/spi/count_s_389\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[0]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => ADLIB_VCC1, S => 
        OPEN, Y => OPEN, FCO => \STAMP_0/spi/count_s_389_FCO\, CC
         => NET_CC_CONFIG925, P => NET_CC_CONFIG923, UB => 
        NET_CC_CONFIG924);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_214\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2]\, 
        IPC => OPEN);
    
    \STAMP_0/spi/count[26]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB12_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[26]\);
    
    \STAMP_0/spi/rx_data[13]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[13]\);
    
    \STAMP_0/PRDATA[29]\ : SLE
      port map(D => \STAMP_0/N_679\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_83\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[29]\);
    
    AFLSDF_INV_12 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_12\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_34_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_84\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_34_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_273\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_33\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[11]\, B => 
        \MemorySynchronizer_0/un104_in_enable_10\, C => 
        \MemorySynchronizer_0/un104_in_enable_11\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[10]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[4]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[5]\, CC
         => NET_CC_CONFIG553, P => NET_CC_CONFIG551, UB => 
        NET_CC_CONFIG552);
    
    \STAMP_0/spi/state[0]\ : SLE
      port map(D => \STAMP_0/spi/busy_7\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/state_Z[0]\);
    
    \MemorySynchronizer_0/ConfigReg[9]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[9]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_21_RNI4G2E8\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[23]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[22]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[23]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[22]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[10]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[11]\, CC
         => NET_CC_CONFIG1150, P => NET_CC_CONFIG1148, UB => 
        NET_CC_CONFIG1149);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_18\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[27]\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[17]\, C => 
        \MemorySynchronizer_0/waitingtimercounter_Z[9]\, D => 
        \MemorySynchronizer_0/waitingtimercounter_Z[3]\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_18_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \MemorySynchronizer_0/TimeStampValue[0]\, Y
         => \MemorySynchronizer_0/TimeStampGen/counter_s[0]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_137\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_35_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[30]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_35_i\);
    
    \STAMP_0/spi/un7_count_NE_18\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \STAMP_0/spi/count_Z[11]\, B => 
        \STAMP_0/spi/count_Z[10]\, C => \STAMP_0/spi/count_Z[9]\, 
        D => \STAMP_0/spi/count_Z[8]\, Y => 
        \STAMP_0/spi/un7_count_NE_18_Z\);
    
    \STAMP_0/spi/count_cry[13]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[13]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[12]\, S => 
        \STAMP_0/spi/count_s[13]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[13]\, CC => NET_CC_CONFIG964, P
         => NET_CC_CONFIG962, UB => NET_CC_CONFIG963);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_82\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/TimeStampGen/prescaler[2]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc2_Z\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[2]\);
    
    \STAMP_0/delay_counter_lm_0[0]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/delay_counter_cry_Y[0]\, B => 
        \STAMP_0/apb_spi_finished_0_sqmuxa_1\, C => 
        \STAMP_0/component_state_RNIFR114_Z[0]\, Y => 
        \STAMP_0/delay_counter_lm[0]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[20]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[20]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[22]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[20]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_61_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_85\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_61_set_Z\);
    
    \STAMP_0/un5_async_prescaler_count_cry_4\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[4]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_3_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_4_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_4_Z\, CC
         => NET_CC_CONFIG492, P => NET_CC_CONFIG490, UB => 
        NET_CC_CONFIG491);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_207\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/SynchStatusReg[29]\ : SLE
      port map(D => \MemorySynchronizer_0/N_113_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[29]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[1]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[1]\);
    
    \MemorySynchronizer_0/SynchStatusReg_152s2_0_0\ : CFG4
      generic map(INIT => x"AFBF")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[2]\, 
        B => \MemorySynchronizer_0/MemorySyncState_Z[0]\, C => 
        ENABLE_MEMORY_LED_c, D => 
        \MemorySynchronizer_0/MemorySyncState_Z[1]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_152_sm0\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_172\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_45_FCINST1\ : 
        FCEND_BUFF_CC
      port map(FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_I_45_FCNET1\, CO
         => \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, 
        CC => NET_CC_CONFIG586, P => NET_CC_CONFIG584, UB => 
        NET_CC_CONFIG585);
    
    \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_0\ : 
        CFG4
      generic map(INIT => x"CD05")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => \MemorySynchronizer_0/APBState_Z[0]\, C => 
        \MemorySynchronizer_0/un1_enabletimestampgen2_2_sn\, D
         => \MemorySynchronizer_0/N_2594\, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_0_Z\);
    
    \STAMP_0/un1_spi_rx_data_0[17]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[17]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[17]\, Y
         => \STAMP_0/N_600\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_11\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[11]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_10_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[21]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_11_Z\, CC
         => NET_CC_CONFIG330, P => NET_CC_CONFIG328, UB => 
        NET_CC_CONFIG329);
    
    \MemorySynchronizer_0/un104_in_enable_cry_11\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[11]\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[11]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_10_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_11_Z\, CC => 
        NET_CC_CONFIG856, P => NET_CC_CONFIG854, UB => 
        NET_CC_CONFIG855);
    
    \MMUART_0_TXD_M2F_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => MMUART_0_TXD_M2F, D => 
        \MMUART_0_TXD_M2F_obuf/U0/DOUT\, E => 
        \MMUART_0_TXD_M2F_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_56_set_RNIPQVF\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_56_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[6]\, C => 
        \MemorySynchronizer_0/un1_nreset_49_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[6]\);
    
    \STAMP_0/spi/count_lm_0[9]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[9]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[9]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[21]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[21]\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_0_CC_2\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO624, CO => OPEN, P(0) => 
        NET_CC_CONFIG694, P(1) => NET_CC_CONFIG697, P(2) => 
        NET_CC_CONFIG700, P(3) => NET_CC_CONFIG703, P(4) => 
        NET_CC_CONFIG706, P(5) => NET_CC_CONFIG709, P(6) => 
        NET_CC_CONFIG712, P(7) => NET_CC_CONFIG715, P(8) => 
        NET_CC_CONFIG718, P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, 
        P(11) => ADLIB_VCC1, UB(0) => NET_CC_CONFIG695, UB(1) => 
        NET_CC_CONFIG698, UB(2) => NET_CC_CONFIG701, UB(3) => 
        NET_CC_CONFIG704, UB(4) => NET_CC_CONFIG707, UB(5) => 
        NET_CC_CONFIG710, UB(6) => NET_CC_CONFIG713, UB(7) => 
        NET_CC_CONFIG716, UB(8) => NET_CC_CONFIG719, UB(9) => 
        ADLIB_VCC1, UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, 
        CC(0) => NET_CC_CONFIG696, CC(1) => NET_CC_CONFIG699, 
        CC(2) => NET_CC_CONFIG702, CC(3) => NET_CC_CONFIG705, 
        CC(4) => NET_CC_CONFIG708, CC(5) => NET_CC_CONFIG711, 
        CC(6) => NET_CC_CONFIG714, CC(7) => NET_CC_CONFIG717, 
        CC(8) => NET_CC_CONFIG720, CC(9) => nc394, CC(10) => nc32, 
        CC(11) => nc40);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13[28]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_0_Z[28]\, B
         => \MemorySynchronizer_0/N_271\, C => 
        \sb_sb_0_STAMP_PADDR[3]\, D => \sb_sb_0_STAMP_PADDR[6]\, 
        Y => \MemorySynchronizer_0/N_2595\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_275\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PRESET_N_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter[11]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[11]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_55_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[11]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_23\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un104_in_enable_23\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[23]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_22_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_23_Z\, CC => 
        NET_CC_CONFIG892, P => NET_CC_CONFIG890, UB => 
        NET_CC_CONFIG891);
    
    \STAMP_0/status_temp_overwrittenVal\ : SLE
      port map(D => \STAMP_0/status_temp_overwrittenVal_9_Z\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN
         => \STAMP_0/un1_new_avail_0_sqmuxa_2_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[10]\);
    
    \STAMP_0/delay_counter_RNI2HNK2[10]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \STAMP_0/N_517_i_0_a2_19\, B => 
        \STAMP_0/N_517_i_0_a2_18\, C => \STAMP_0/N_517_i_0_a2_17\, 
        D => \STAMP_0/N_517_i_0_a2_16\, Y => 
        \STAMP_0/N_517_i_0_a2_25\);
    
    \MemorySynchronizer_0/TimeStampReg[23]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[23]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[23]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[17]\ : SLE
      port map(D => \STAMP_0_data_frame[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[17]\);
    
    \STAMP_0/spi/count_cry[2]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[2]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[1]\, S => 
        \STAMP_0/spi/count_s[2]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[2]\, CC => NET_CC_CONFIG931, P
         => NET_CC_CONFIG929, UB => NET_CC_CONFIG930);
    
    \MemorySynchronizer_0/un94_in_enable_28\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/un94_in_enable_19_Z\, B
         => \MemorySynchronizer_0/un94_in_enable_18_Z\, C => 
        \MemorySynchronizer_0/un94_in_enable_17_Z\, D => 
        \MemorySynchronizer_0/un94_in_enable_16_Z\, Y => 
        \MemorySynchronizer_0/un94_in_enable_28_Z\);
    
    \STAMP_0/spi/tx_buffer[1]\ : SLE
      port map(D => \STAMP_0/spi/N_140\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[1]\);
    
    \MemorySynchronizer_0/un94_in_enable_17\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[22]\, B => 
        \MemorySynchronizer_0/resettimercounter_Z[21]\, C => 
        \MemorySynchronizer_0/resettimercounter_Z[20]\, D => 
        \MemorySynchronizer_0/resettimercounter_Z[19]\, Y => 
        \MemorySynchronizer_0/un94_in_enable_17_Z\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[6]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[6]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[30]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_30_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[2]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_CC_2\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO101, CO => OPEN, P(0) => 
        NET_CC_CONFIG171, P(1) => NET_CC_CONFIG174, P(2) => 
        NET_CC_CONFIG177, P(3) => NET_CC_CONFIG180, P(4) => 
        NET_CC_CONFIG183, P(5) => NET_CC_CONFIG186, P(6) => 
        NET_CC_CONFIG189, P(7) => NET_CC_CONFIG192, P(8) => 
        ADLIB_VCC1, P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, 
        P(11) => ADLIB_VCC1, UB(0) => NET_CC_CONFIG172, UB(1) => 
        NET_CC_CONFIG175, UB(2) => NET_CC_CONFIG178, UB(3) => 
        NET_CC_CONFIG181, UB(4) => NET_CC_CONFIG184, UB(5) => 
        NET_CC_CONFIG187, UB(6) => NET_CC_CONFIG190, UB(7) => 
        NET_CC_CONFIG193, UB(8) => ADLIB_VCC1, UB(9) => 
        ADLIB_VCC1, UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, 
        CC(0) => NET_CC_CONFIG173, CC(1) => NET_CC_CONFIG176, 
        CC(2) => NET_CC_CONFIG179, CC(3) => NET_CC_CONFIG182, 
        CC(4) => NET_CC_CONFIG185, CC(5) => NET_CC_CONFIG188, 
        CC(6) => NET_CC_CONFIG191, CC(7) => NET_CC_CONFIG194, 
        CC(8) => nc297, CC(9) => nc99, CC(10) => nc75, CC(11) => 
        nc183);
    
    \STAMP_0/un1_spi_rx_data[6]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_656\, C => \STAMP_0/spi_rx_data[6]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[6]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_108\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0]\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/spi/count[23]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[23]\);
    
    \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1_0_a2_1\ : 
        CFG3
      generic map(INIT => x"EF")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, C => \sb_sb_0_STAMP_PADDR[4]\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1_0_a2_1_Z\);
    
    \STAMP_0/un1_spi_rx_data_2[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_588\, B => \STAMP_0/N_622\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_655\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_184\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net\, 
        IPC => OPEN);
    
    AFLSDF_INV_35 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_35\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_1_1[4]\ : 
        CFG4
      generic map(INIT => x"4000")

      port map(A => STAMP_0_new_avail, B => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_28_Z\, 
        C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_29_Z\, 
        D => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, Y
         => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_1_1_Z[4]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[17]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[17]\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/N_2323\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[17]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[17]\);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB3\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[13]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => \MemorySynchronizer_0/N_2597\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[13]\, C => 
        \MemorySynchronizer_0/TimeStampReg_Z[13]\, D => 
        \MemorySynchronizer_0/N_1236\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[13]\);
    
    \MemorySynchronizer_0/un94_in_enable_21\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[8]\, 
        B => \MemorySynchronizer_0/resettimercounter_Z[7]\, C => 
        \MemorySynchronizer_0/resettimercounter_Z[6]\, D => 
        \MemorySynchronizer_0/resettimercounter_Z[5]\, Y => 
        \MemorySynchronizer_0/un94_in_enable_21_Z\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_23\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[26]\, B => 
        \MemorySynchronizer_0/un120_in_enable_i_A[27]\, C => 
        \MemorySynchronizer_0/un120_in_enable_i_A[28]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[29]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_23_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[20]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[20]\, B => 
        \MemorySynchronizer_0/un104_in_enable_20\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[20]\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_YR\);
    
    \MemorySynchronizer_0/SynchStatusReg2[13]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[13]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[13]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_243\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3]\, IPC
         => OPEN);
    
    \STAMP_0/delay_counter_cry[2]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[2]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/delay_counter_cry_Z[1]\, S => 
        \STAMP_0/delay_counter_s[2]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[2]\, CC => NET_CC_CONFIG401, 
        P => NET_CC_CONFIG399, UB => NET_CC_CONFIG400);
    
    \STAMP_0/dummy[20]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_86\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[20]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[21]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[21]\, B => 
        \sb_sb_0_STAMP_PWDATA[21]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[21]\);
    
    \MemorySynchronizer_0/un1_nreset_17_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_44_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_17_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_17_rs_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_85\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[1]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[20]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[20]\, B => 
        \sb_sb_0_STAMP_PWDATA[20]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[20]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[0]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[0]\, B => 
        \MemorySynchronizer_0/un104_in_enable_0\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[0]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_59\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20]\, 
        IPC => OPEN);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[27]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[27]\, B => 
        \sb_sb_0_Memory_PRDATA[27]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[27]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_210\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter_0_sqmuxa_1_0_a2\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, B => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, C => 
        ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/resettimercounter_0_sqmuxa_1\);
    
    \MemorySynchronizer_0/un1_nreset_11_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_38_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_11_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_11_rs_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[1]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[1]\, B => 
        \MemorySynchronizer_0/un104_in_enable_1\, C => 
        \MemorySynchronizer_0/N_2574\, D => 
        \MemorySynchronizer_0/N_2577\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[1]\);
    
    \STAMP_0/async_prescaler_count[0]\ : SLE
      port map(D => \STAMP_0/async_prescaler_count_5_Z[0]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => \AND2_0_RNIKOS1/U0_RGB1_YR\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/async_prescaler_count_Z[0]\);
    
    \MemorySynchronizer_0/TimeStampReg[13]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[13]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[13]\);
    
    \STAMP_0/un1_spi_rx_data_2[11]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_594\, B => \STAMP_0/N_628\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_661\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_79\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20]\, 
        IPC => OPEN);
    
    \RXSM_SOE_ibuf/U0/U_IOINFF\ : IOINFF_BYPASS
      port map(A => \RXSM_SOE_ibuf/U0/YIN1\, Y => 
        \RXSM_SOE_ibuf/U0/YIN\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[16]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_16_S\, 
        Y => \MemorySynchronizer_0/N_1517\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1[2]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => \MemorySynchronizer_0/N_2510\, B => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_0_0_0[4]\, 
        C => \MemorySynchronizer_0/SynchStatusReg_Z[4]\, D => 
        \MemorySynchronizer_0/N_2606\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168[2]\);
    
    \STAMP_0/config[18]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[18]\);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[0]\ : 
        CFG2
      generic map(INIT => x"6")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[0]\, Y => 
        \MemorySynchronizer_0/N_1091\);
    
    \MemorySynchronizer_0/SynchStatusReg2[26]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_RNO_Z[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[26]\);
    
    \MemorySynchronizer_0/un1_nreset_25_rs_RNI2LG6\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_37_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[23]\, C
         => \MemorySynchronizer_0/un1_nreset_25_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[23]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[1]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_1_S\, 
        Y => \MemorySynchronizer_0/N_1561\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[17]\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \MemorySynchronizer_0/N_2577\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[17]\, C => 
        \MemorySynchronizer_0/un104_in_enable_17\, D => 
        \MemorySynchronizer_0/N_1445\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[17]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_19\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[19]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[19]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_18\, S => 
        \MemorySynchronizer_0/temp_1[19]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_19\, CC => 
        NET_CC_CONFIG256, P => NET_CC_CONFIG254, UB => 
        NET_CC_CONFIG255);
    
    \nCS2_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \nCS2_obuf/U0/DOUT1\, Y => 
        \nCS2_obuf/U0/DOUT\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_0_CC_0\ : 
        CC_CONFIG
      port map(CI => ADLIB_GND0, CO => CI_TO_CO721, P(0) => 
        NET_CC_CONFIG723, P(1) => NET_CC_CONFIG726, P(2) => 
        NET_CC_CONFIG729, P(3) => NET_CC_CONFIG732, P(4) => 
        NET_CC_CONFIG735, P(5) => NET_CC_CONFIG738, P(6) => 
        NET_CC_CONFIG741, P(7) => NET_CC_CONFIG744, P(8) => 
        NET_CC_CONFIG747, P(9) => NET_CC_CONFIG750, P(10) => 
        NET_CC_CONFIG753, P(11) => NET_CC_CONFIG756, UB(0) => 
        NET_CC_CONFIG724, UB(1) => NET_CC_CONFIG727, UB(2) => 
        NET_CC_CONFIG730, UB(3) => NET_CC_CONFIG733, UB(4) => 
        NET_CC_CONFIG736, UB(5) => NET_CC_CONFIG739, UB(6) => 
        NET_CC_CONFIG742, UB(7) => NET_CC_CONFIG745, UB(8) => 
        NET_CC_CONFIG748, UB(9) => NET_CC_CONFIG751, UB(10) => 
        NET_CC_CONFIG754, UB(11) => NET_CC_CONFIG757, CC(0) => 
        NET_CC_CONFIG725, CC(1) => NET_CC_CONFIG728, CC(2) => 
        NET_CC_CONFIG731, CC(3) => NET_CC_CONFIG734, CC(4) => 
        NET_CC_CONFIG737, CC(5) => NET_CC_CONFIG740, CC(6) => 
        NET_CC_CONFIG743, CC(7) => NET_CC_CONFIG746, CC(8) => 
        NET_CC_CONFIG749, CC(9) => NET_CC_CONFIG752, CC(10) => 
        NET_CC_CONFIG755, CC(11) => NET_CC_CONFIG758);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[5]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[5]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_142\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net\, IPC
         => OPEN);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_49_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[1]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_49\);
    
    \MemorySynchronizer_0/SynchStatusReg[22]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_34_Z[20]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[22]\);
    
    \MemorySynchronizer_0/un1_nreset_2_rs_RNITBF11\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_48_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[3]\, C
         => \MemorySynchronizer_0/un1_nreset_2_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[3]\);
    
    \debug_led_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \debug_led_obuf/U0/EOUT1\, Y => 
        \debug_led_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv[27]\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_27\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[27]\, 
        C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[4]\, D
         => \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, 
        Y => \MemorySynchronizer_0/waitingtimercounter_10[27]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[18]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[18]\, B => 
        \sb_sb_0_STAMP_PWDATA[18]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[18]\);
    
    AFLSDF_INV_74 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_74\);
    
    \STAMP_0/un1_spi_rx_data_2[0]\ : CFG4
      generic map(INIT => x"D155")

      port map(A => \STAMP_0/un1_spi_rx_data_2_1_0_Z[0]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/dummy_Z[0]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_650\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[6]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[6]\);
    
    \STAMP_0/status_temp_newVal\ : SLE
      port map(D => \STAMP_0/drdy_flank_detected_temp_1_sqmuxa_1\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \STAMP_0/un1_new_avail_0_sqmuxa_2_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[13]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[19]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[19]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[19]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[19]\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_15\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[15]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_14_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[17]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_15_Z\, CC
         => NET_CC_CONFIG342, P => NET_CC_CONFIG340, UB => 
        NET_CC_CONFIG341);
    
    \MemorySynchronizer_0/ConfigReg[7]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[7]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_35\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[14]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_35_Z\);
    
    
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_29\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_20_Z\, 
        B => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_23_Z\, 
        C => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_22_Z\, 
        D => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_21_Z\, 
        Y => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_29_Z\);
    
    \STAMP_0/spi/mosi_1_1_0_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/mosi_1_1_2\, B => 
        debug_led_net_0, C => \STAMP_0/spi/un10_count_i\, Y => 
        \STAMP_0/spi/mosi_1_1\);
    
    \STAMP_0/measurement_dms2[7]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[39]\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\);
    
    \STAMP_0/spi/count_cry[11]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[11]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[10]\, S => 
        \STAMP_0/spi/count_s[11]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[11]\, CC => NET_CC_CONFIG958, P
         => NET_CC_CONFIG956, UB => NET_CC_CONFIG957);
    
    \STAMP_0/un1_apb_spi_finished_1_f0\ : CFG3
      generic map(INIT => x"54")

      port map(A => \STAMP_0/apb_spi_finished_0_sqmuxa\, B => 
        \STAMP_0/apb_spi_finished_Z\, C => 
        \STAMP_0/apb_spi_finished_1_sqmuxa\, Y => 
        \STAMP_0/un1_apb_spi_finished_1_f0_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_245\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5]\, IPC
         => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_RNO[27]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_27_S\, 
        Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[4]\);
    
    \STAMP_0/delay_counter_lm_0[22]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[22]\, Y => 
        \STAMP_0/delay_counter_lm[22]\);
    
    \MemorySynchronizer_0/PRDATA[4]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[4]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[27]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[27]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[27]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[26]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_26\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_208\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0[28]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/N_1168\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[28]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[28]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[28]\, Y => 
        \MemorySynchronizer_0/PRDATA_21[28]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_17\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[22]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[29]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[28]\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[28]\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[28]\, C => 
        \MemorySynchronizer_0/N_2593\, D => 
        \MemorySynchronizer_0/N_1163\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[28]\);
    
    \adc_clk_obuf/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \adc_clk_obuf/U0/EOUT1\, Y => 
        \adc_clk_obuf/U0/EOUT\);
    
    \STAMP_0/spi/count_s_389_CC_2\ : CC_CONFIG
      port map(CI => CI_TO_CO921, CO => CI_TO_CO922, P(0) => 
        NET_CC_CONFIG962, P(1) => NET_CC_CONFIG965, P(2) => 
        NET_CC_CONFIG968, P(3) => NET_CC_CONFIG971, P(4) => 
        NET_CC_CONFIG974, P(5) => NET_CC_CONFIG977, P(6) => 
        NET_CC_CONFIG980, P(7) => NET_CC_CONFIG983, P(8) => 
        NET_CC_CONFIG986, P(9) => NET_CC_CONFIG989, P(10) => 
        NET_CC_CONFIG992, P(11) => NET_CC_CONFIG995, UB(0) => 
        NET_CC_CONFIG963, UB(1) => NET_CC_CONFIG966, UB(2) => 
        NET_CC_CONFIG969, UB(3) => NET_CC_CONFIG972, UB(4) => 
        NET_CC_CONFIG975, UB(5) => NET_CC_CONFIG978, UB(6) => 
        NET_CC_CONFIG981, UB(7) => NET_CC_CONFIG984, UB(8) => 
        NET_CC_CONFIG987, UB(9) => NET_CC_CONFIG990, UB(10) => 
        NET_CC_CONFIG993, UB(11) => NET_CC_CONFIG996, CC(0) => 
        NET_CC_CONFIG964, CC(1) => NET_CC_CONFIG967, CC(2) => 
        NET_CC_CONFIG970, CC(3) => NET_CC_CONFIG973, CC(4) => 
        NET_CC_CONFIG976, CC(5) => NET_CC_CONFIG979, CC(6) => 
        NET_CC_CONFIG982, CC(7) => NET_CC_CONFIG985, CC(8) => 
        NET_CC_CONFIG988, CC(9) => NET_CC_CONFIG991, CC(10) => 
        NET_CC_CONFIG994, CC(11) => NET_CC_CONFIG997);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[22]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[22]\, B => 
        \sb_sb_0_Memory_PRDATA[22]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[22]\);
    
    \MemorySynchronizer_0/PRDATA[22]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[22]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[22]\);
    
    \MemorySynchronizer_0/un105_in_enable_i_0_a2_15\ : CFG3
      generic map(INIT => x"01")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[30]\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[10]\, C => 
        \MemorySynchronizer_0/waitingtimercounter_Z[0]\, Y => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_15_Z\);
    
    \MemorySynchronizer_0/un1_nreset_37_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_44\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_37_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_37_rs_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[24]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[24]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[24]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[10]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \MemorySynchronizer_0/N_2585\, B => 
        \MemorySynchronizer_0/N_2581\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[10]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[10]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0[10]\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_9\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[3]\, 
        B => \MemorySynchronizer_0/un104_in_enable_2\, C => 
        \MemorySynchronizer_0/un104_in_enable_3\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[2]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[0]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[1]\, CC
         => NET_CC_CONFIG541, P => NET_CC_CONFIG539, UB => 
        NET_CC_CONFIG540);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[12]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[12]\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2564\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1469\);
    
    \STAMP_0/spi/rx_buffer[11]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[11]\);
    
    \MemorySynchronizer_0/waitingtimercounter[7]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_59_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[7]\);
    
    \MemorySynchronizer_0/un1_nreset_31_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/N_1978_i\, EN => ADLIB_VCC1, ALn
         => \MemorySynchronizer_0/un1_nreset_31_i\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_31_rs_Z\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_7\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/CLK3_net\, IPB => OPEN, 
        IPC => \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[5]\);
    
    \MemorySynchronizer_0/TimeStampReg[26]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[26]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[26]\);
    
    \STAMP_0/delay_counter_cry[20]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[20]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[19]\, S
         => \STAMP_0/delay_counter_s[20]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[20]\, CC => NET_CC_CONFIG455, 
        P => NET_CC_CONFIG453, UB => NET_CC_CONFIG454);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[23]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[23]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[22]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[23]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[23]\, CC
         => NET_CC_CONFIG75, P => NET_CC_CONFIG73, UB => 
        NET_CC_CONFIG74);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_a2_0[1]\ : 
        CFG2
      generic map(INIT => x"4")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, B => 
        \MemorySynchronizer_0/SynchStatusReg_Z[3]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_a2_0_Z[1]\);
    
    AFLSDF_INV_99 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_54_i_i_a2_Z\, 
        Y => \AFLSDF_INV_99\);
    
    \MemorySynchronizer_0/un1_nreset_53_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[13]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_53_i\);
    
    \STAMP_0/un1_spi_rx_data_2[23]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_606\, B => \STAMP_0/N_640\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_673\);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB1\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB1_rgbr_net_1\);
    
    AFLSDF_INV_42 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_40\, Y => 
        \AFLSDF_INV_42\);
    
    \STAMP_0/component_state_ns_0_i_0_tz[0]\ : CFG4
      generic map(INIT => x"880F")

      port map(A => \STAMP_0/spi_request_for_Z[0]\, B => 
        \STAMP_0/spi_request_for_Z[1]\, C => 
        \STAMP_0/component_state_Z[5]\, D => 
        \STAMP_0/component_state_Z[0]\, Y => 
        \STAMP_0/component_state_ns_0_i_0_tz_Z[0]\);
    
    AFLSDF_INV_97 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_50\, Y => 
        \AFLSDF_INV_97\);
    
    \MOSI_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => MOSI_c, E => ADLIB_VCC1, DOUT => 
        \MOSI_obuf/U0/DOUT1\, EOUT => \MOSI_obuf/U0/EOUT1\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_35_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_87\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_35_set_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[12]\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \MemorySynchronizer_0/N_2577\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[12]\, C => 
        \MemorySynchronizer_0/un104_in_enable_12\, D => 
        \MemorySynchronizer_0/N_1469\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[12]\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_75\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[9]\, 
        B => \MemorySynchronizer_0/un104_in_enable_8\, C => 
        \MemorySynchronizer_0/un104_in_enable_9\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[8]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[3]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[4]\, CC
         => NET_CC_CONFIG550, P => NET_CC_CONFIG548, UB => 
        NET_CC_CONFIG549);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[7]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[1]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[7]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[7]\);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB5\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[25]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[25]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[25]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[25]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_171\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_17_RNI7UO58\ : 
        ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[19]\, B => 
        \MemorySynchronizer_0/un120_in_enable_a_4[18]\, C => 
        \MemorySynchronizer_0/un120_in_enable_a_4[19]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[18]\, FCI => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[8]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[9]\, CC
         => NET_CC_CONFIG1144, P => NET_CC_CONFIG1142, UB => 
        NET_CC_CONFIG1143);
    
    \STAMP_0/async_state[1]\ : SLE
      port map(D => \STAMP_0/async_state_17[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/async_state_Z[1]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_14\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[14]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[14]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_13\, S => 
        \MemorySynchronizer_0/temp_1[14]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_14\, CC => 
        NET_CC_CONFIG241, P => NET_CC_CONFIG239, UB => 
        NET_CC_CONFIG240);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[12]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[12]\);
    
    \STAMP_0/status_async_cycles_lm_0[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/status_async_cycles_3_sqmuxa\, B => 
        \STAMP_0/status_async_cycles_s[4]\, C => 
        \STAMP_0/status_async_cycles_1_sqmuxa_Z\, Y => 
        \STAMP_0/status_async_cycles_lm[4]\);
    
    \MemorySynchronizer_0/waitingtimercounter[28]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[28]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_37_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[28]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[31]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s_Z[31]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[31]\);
    
    \STAMP_0/delay_counter_cry[7]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => \STAMP_0/delay_counter_Z[7]\, 
        C => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/delay_counter_cry_Z[6]\, S => 
        \STAMP_0/delay_counter_s[7]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[7]\, CC => NET_CC_CONFIG416, 
        P => NET_CC_CONFIG414, UB => NET_CC_CONFIG415);
    
    \STAMP_0/async_prescaler_count_5[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \STAMP_0/un1_async_prescaler_count\, B => 
        \STAMP_0/un5_async_prescaler_count_cry_8_S\, Y => 
        \STAMP_0/async_prescaler_count_5_Z[8]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_226\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/TimeStampGen/prescaler[3]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_5_Z[3]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[3]\);
    
    \STAMP_0/spi/clk_toggles_lm_0[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/spi/ss_n_buffer_1_sqmuxa\, B => 
        \STAMP_0/spi/clk_toggles_s[4]\, Y => 
        \STAMP_0/spi/clk_toggles_lm[4]\);
    
    \MemorySynchronizer_0/un1_nreset_55_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_55\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_55_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_55_rs_Z\);
    
    \MemorySynchronizer_0/ConfigReg[27]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[27]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[27]\);
    
    \MemorySynchronizer_0/resynctimercounter[8]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1114\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[8]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[2]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_2_S\, 
        Y => \MemorySynchronizer_0/N_1565\);
    
    \MemorySynchronizer_0/resynctimercounter[24]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1098\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[24]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_27\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_19\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_12_S\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_13_S\, 
        C => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_14_S\, D
         => \MemorySynchronizer_0/un5_resettimercounter_cry_15_S\, 
        Y => \MemorySynchronizer_0/un6_in_enable_0_a3_19_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_RNO[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[6]\, Y => 
        \MemorySynchronizer_0/ResetTimerValueReg_m_0_0[6]\);
    
    AFLSDF_INV_31 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_31\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[4]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[4]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[3]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[4]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[4]\, CC
         => NET_CC_CONFIG18, P => NET_CC_CONFIG16, UB => 
        NET_CC_CONFIG17);
    
    \MemorySynchronizer_0/un104_in_enable_cry_31_RNISAUC\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/un104_in_enable_cry_31_Z\, B => 
        \MemorySynchronizer_0/un104_in_enable_axb_31\, Y => 
        \MemorySynchronizer_0/un105_m1_e_0_0\);
    
    \MemorySynchronizer_0/numberofnewavails_RNIVL541_1[0]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[2]\, 
        B => \MemorySynchronizer_0/numberofnewavails_Z[1]\, C => 
        \MemorySynchronizer_0/numberofnewavails_Z[0]\, Y => 
        \MemorySynchronizer_0/numberofnewavails_RNIVL541_1_Z[0]\);
    
    \MemorySynchronizer_0/TimeStampReg[16]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[16]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[16]\);
    
    \MemorySynchronizer_0/numberofpendingresyncrequest[1]\ : SLE
      port map(D => \MemorySynchronizer_0/ConfigReg_Z[5]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN
         => \MemorySynchronizer_0/numberofnewavails_0_sqmuxa\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/numberofpendingresyncrequest_Z[1]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_2[20]\ : 
        CFG2
      generic map(INIT => x"1")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[2]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[4]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_2_Z[20]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_217\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25]\);
    
    \MemorySynchronizer_0/waitingtimercounter[2]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_45_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[2]\);
    
    \STAMP_0/delay_counter_lm_0[16]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[16]\, Y => 
        \STAMP_0/delay_counter_lm[16]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_222\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_14\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[19]\, B
         => ADLIB_VCC1, C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19]\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/delay_counter_cry[19]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[19]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[18]\, S
         => \STAMP_0/delay_counter_s[19]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[19]\, CC => NET_CC_CONFIG452, 
        P => NET_CC_CONFIG450, UB => NET_CC_CONFIG451);
    
    \MemorySynchronizer_0/ConfigReg[14]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[14]\);
    
    \STAMP_0/measurement_temp[7]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[23]\);
    
    \MemorySynchronizer_0/resettimercounter[25]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_29_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[25]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[4]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_4_S\, 
        Y => \MemorySynchronizer_0/N_1549\);
    
    \STAMP_0/delay_counter[13]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[13]\);
    
    \stamp0_spi_temp_cs_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => stamp0_spi_temp_cs_c, E => ADLIB_VCC1, DOUT
         => \stamp0_spi_temp_cs_obuf/U0/DOUT1\, EOUT => 
        \stamp0_spi_temp_cs_obuf/U0/EOUT1\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[19]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[19]\);
    
    \STAMP_0/spi/count_cry[6]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[6]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[5]\, S => 
        \STAMP_0/spi/count_s[6]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[6]\, CC => NET_CC_CONFIG943, P
         => NET_CC_CONFIG941, UB => NET_CC_CONFIG942);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_0_CC_2\ : 
        CC_CONFIG
      port map(CI => CI_TO_CO196, CO => OPEN, P(0) => 
        NET_CC_CONFIG263, P(1) => NET_CC_CONFIG266, P(2) => 
        NET_CC_CONFIG269, P(3) => NET_CC_CONFIG272, P(4) => 
        NET_CC_CONFIG275, P(5) => NET_CC_CONFIG278, P(6) => 
        NET_CC_CONFIG281, P(7) => NET_CC_CONFIG284, P(8) => 
        NET_CC_CONFIG287, P(9) => NET_CC_CONFIG290, P(10) => 
        ADLIB_VCC1, P(11) => ADLIB_VCC1, UB(0) => 
        NET_CC_CONFIG264, UB(1) => NET_CC_CONFIG267, UB(2) => 
        NET_CC_CONFIG270, UB(3) => NET_CC_CONFIG273, UB(4) => 
        NET_CC_CONFIG276, UB(5) => NET_CC_CONFIG279, UB(6) => 
        NET_CC_CONFIG282, UB(7) => NET_CC_CONFIG285, UB(8) => 
        NET_CC_CONFIG288, UB(9) => NET_CC_CONFIG291, UB(10) => 
        ADLIB_VCC1, UB(11) => ADLIB_VCC1, CC(0) => 
        NET_CC_CONFIG265, CC(1) => NET_CC_CONFIG268, CC(2) => 
        NET_CC_CONFIG271, CC(3) => NET_CC_CONFIG274, CC(4) => 
        NET_CC_CONFIG277, CC(5) => NET_CC_CONFIG280, CC(6) => 
        NET_CC_CONFIG283, CC(7) => NET_CC_CONFIG286, CC(8) => 
        NET_CC_CONFIG289, CC(9) => NET_CC_CONFIG292, CC(10) => 
        nc435, CC(11) => nc345);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[14]\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \MemorySynchronizer_0/N_2577\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[14]\, C => 
        \MemorySynchronizer_0/un104_in_enable_14\, D => 
        \MemorySynchronizer_0/N_1461\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[14]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[7]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_64\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[7]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[7]\, D
         => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[7]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/N_2564\, B => 
        \MemorySynchronizer_0/N_2561\, C => 
        \MemorySynchronizer_0/APBState_Z[1]\, D => 
        \sb_sb_0_STAMP_PADDR[6]\, Y => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\);
    
    \MemorySynchronizer_0/un1_nreset_40_rs_RNIUP7G\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_31_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[19]\, C
         => \MemorySynchronizer_0/un1_nreset_40_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[19]\);
    
    \STAMP_0/spi/rx_buffer[14]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[14]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_55\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[27]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_55_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[22]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[22]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[24]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[22]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[26]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[26]\, B => 
        \sb_sb_0_STAMP_PWDATA[26]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[26]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_17\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_18\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_16_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[18]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_17_Z\, CC
         => NET_CC_CONFIG1074, P => NET_CC_CONFIG1072, UB => 
        NET_CC_CONFIG1073);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[7]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[7]\, C => 
        \MemorySynchronizer_0/resynctimercounter_1[25]\, Y => 
        \MemorySynchronizer_0/N_1084\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_12[17]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[17]\, B => 
        \sb_sb_0_STAMP_PADDR[6]\, C => 
        \MemorySynchronizer_0/N_2564\, D => 
        \MemorySynchronizer_0/N_2561\, Y => 
        \MemorySynchronizer_0/N_1445\);
    
    \STAMP_0/un1_spi_rx_data_1[21]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[53]\, B => 
        \STAMP_0/dummy_Z[21]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_638\);
    
    \MemorySynchronizer_0/resynctimercounter[20]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1102\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[20]\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_3_0[20]\ : 
        CFG3
      generic map(INIT => x"0E")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\, 
        C => \MemorySynchronizer_0/SynchStatusReg_Z[25]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_3_0_Z[20]\);
    
    \MemorySynchronizer_0/N_2533_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_88\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_2533_set_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc5\ : 
        CFG3
      generic map(INIT => x"78")

      port map(A => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[4]\, B => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_c4\, C
         => \MemorySynchronizer_0/TimeStampGen/prescaler_Z[5]\, Y
         => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc5_Z\);
    
    \STAMP_0/spi/count_lm_0[23]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[23]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[23]\);
    
    \MemorySynchronizer_0/resettimercounter_RNIH6GE[5]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_57_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[5]\, C => 
        \MemorySynchronizer_0/un1_nreset_50_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[5]\);
    
    \MemorySynchronizer_0/resettimercounter_RNIL18V[20]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_40_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[20]\, C => 
        \MemorySynchronizer_0/un1_nreset_13_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[20]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[19]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[19]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_279\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_118\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7]\, 
        IPC => OPEN);
    
    \STAMP_0/un27_paddr_1\ : CFG4
      generic map(INIT => x"7530")

      port map(A => stamp0_ready_dms2_c, B => stamp0_ready_temp_c, 
        C => \sb_sb_0_STAMP_PADDR[6]\, D => 
        \sb_sb_0_STAMP_PADDR[5]\, Y => \STAMP_0/un27_paddr_1_Z\);
    
    \STAMP_0/un1_spi_rx_data_1[31]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[63]\, B => 
        \STAMP_0/dummy_Z[31]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_648\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_141\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2HCALIB_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net\, IPC
         => OPEN);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_5\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[5]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_4_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[27]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_5_Z\, CC
         => NET_CC_CONFIG312, P => NET_CC_CONFIG310, UB => 
        NET_CC_CONFIG311);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[27]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[27]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[27]\, C => 
        \MemorySynchronizer_0/N_2598\, D => 
        \MemorySynchronizer_0/N_2576\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[27]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[23]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[23]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[23]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[23]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_256\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_56_i_i_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[10]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_56_i_i_a2_Z\);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\);
    
    \STAMP_0/un1_spi_rx_data_0[22]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[22]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[22]\, Y
         => \STAMP_0/N_605\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[14]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_14\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[14]\, 
        C => \MemorySynchronizer_0/N_1529\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[14]\);
    
    \MemorySynchronizer_0/resettimercounter[1]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[1]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_33_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[1]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_164\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_28_0_a3_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[26]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_28_i\);
    
    \MemorySynchronizer_0/resettimercounter[31]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[31]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \ResetAND_RNIMHJB/U0_RGB1_YR\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounter_Z[31]\);
    
    \STAMP_0/spi_tx_data_RNO[6]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[6]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_292_i\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_47_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_89\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_47_set_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[18]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[18]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[18]\, C => 
        \MemorySynchronizer_0/N_2598\, D => 
        \MemorySynchronizer_0/N_2576\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[18]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_6\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[6]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_5_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[6]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_6_Z\, 
        CC => NET_CC_CONFIG122, P => NET_CC_CONFIG120, UB => 
        NET_CC_CONFIG121);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_52\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13]\, 
        IPC => OPEN);
    
    \STAMP_0/spi_tx_data_RNO[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[2]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_296_i\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_a3_1[15]\ : 
        CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_15_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => \MemorySynchronizer_0/N_76\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_24\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0]\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_54_i_i_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[9]\, B => NN_1, 
        Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_54_i_i_a2_Z\);
    
    \STAMP_0/un1_spi_rx_data_2[20]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_603\, B => \STAMP_0/N_637\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_670\);
    
    \STAMP_0/spi_tx_data_RNO[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[0]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_298_i\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[17]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[17]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[17]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[15]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[17]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_RNO[13]\ : 
        CFG2
      generic map(INIT => x"8")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[13]\, Y => 
        \MemorySynchronizer_0/ResetTimerValueReg_m_0_0[13]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[14]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_14\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_49_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_90\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_49_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_72\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6]\, 
        IPB => OPEN, IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_252\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_GND0, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0]\);
    
    \STAMP_0/un1_spi_rx_data_1[14]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[46]\, B => 
        \STAMP_0/dummy_Z[14]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_631\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_15\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[5]\, 
        B => \MemorySynchronizer_0/un104_in_enable_4\, C => 
        \MemorySynchronizer_0/un104_in_enable_5\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[4]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[1]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[2]\, CC
         => NET_CC_CONFIG544, P => NET_CC_CONFIG542, UB => 
        NET_CC_CONFIG543);
    
    \sb_sb_0/SYSRESET_POR/INST_SYSRESET_FF_IP\ : SYSRESET_FF
      port map(UDRCAP => OPEN, UDRSH => OPEN, UDRUPD => OPEN, 
        UIREG(7) => nc333, UIREG(6) => nc288, UIREG(5) => nc85, 
        UIREG(4) => nc27, UIREG(3) => nc108, UIREG(2) => nc396, 
        UIREG(1) => nc402, UIREG(0) => nc325, URSTB => OPEN, 
        UDRCK => OPEN, UTDI => OPEN, POWER_ON_RESET_N => 
        sb_sb_0_POWER_ON_RESET_N, FF_TO_START => ff_to_start_net, 
        FF_DONE => OPEN, UTDO => \sb_sb_0/SYSRESET_POR/UTDO_net\, 
        DEVRST_N => DEVRST_N, TDI => ADLIB_VCC1, TMS => 
        ADLIB_VCC1, TCK => ADLIB_VCC1, TRSTB => ADLIB_VCC1, TDO
         => OPEN);
    
    \STAMP_0/spi/clk_toggles_s_390_CC_0\ : CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => OPEN, P(0) => 
        NET_CC_CONFIG605, P(1) => NET_CC_CONFIG608, P(2) => 
        NET_CC_CONFIG611, P(3) => NET_CC_CONFIG614, P(4) => 
        NET_CC_CONFIG617, P(5) => NET_CC_CONFIG620, P(6) => 
        ADLIB_VCC1, P(7) => ADLIB_VCC1, P(8) => ADLIB_VCC1, P(9)
         => ADLIB_VCC1, P(10) => ADLIB_VCC1, P(11) => ADLIB_VCC1, 
        UB(0) => NET_CC_CONFIG606, UB(1) => NET_CC_CONFIG609, 
        UB(2) => NET_CC_CONFIG612, UB(3) => NET_CC_CONFIG615, 
        UB(4) => NET_CC_CONFIG618, UB(5) => NET_CC_CONFIG621, 
        UB(6) => ADLIB_VCC1, UB(7) => ADLIB_VCC1, UB(8) => 
        ADLIB_VCC1, UB(9) => ADLIB_VCC1, UB(10) => ADLIB_VCC1, 
        UB(11) => ADLIB_VCC1, CC(0) => NET_CC_CONFIG607, CC(1)
         => NET_CC_CONFIG610, CC(2) => NET_CC_CONFIG613, CC(3)
         => NET_CC_CONFIG616, CC(4) => NET_CC_CONFIG619, CC(5)
         => NET_CC_CONFIG622, CC(6) => nc16, CC(7) => nc155, 
        CC(8) => nc51, CC(9) => nc301, CC(10) => nc33, CC(11) => 
        nc443);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[1]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[1]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1090\, Y => 
        \MemorySynchronizer_0/N_1121\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[22]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[22]\, B => 
        \MemorySynchronizer_0/un104_in_enable_22\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[22]\);
    
    \stamp0_spi_dms1_cs_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => stamp0_spi_dms1_cs, D => 
        \stamp0_spi_dms1_cs_obuf/U0/DOUT\, E => 
        \stamp0_spi_dms1_cs_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[23]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[23]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[23]\);
    
    \STAMP_0/spi_tx_data[12]\ : SLE
      port map(D => \STAMP_0/un1_pwdata_Z[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[12]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_8\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6[9]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[9]\, B => 
        \MemorySynchronizer_0/un104_in_enable_9\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[9]\);
    
    \MemorySynchronizer_0/un1_nreset_6\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[30]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_6_i\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_26[10]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \sb_sb_0_STAMP_PADDR[5]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, C => 
        \MemorySynchronizer_0/N_271\, D => 
        \MemorySynchronizer_0/N_2567\, Y => 
        \MemorySynchronizer_0/N_2582\);
    
    \STAMP_0/dummy[3]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_91\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[3]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[27]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[27]\, B => 
        \sb_sb_0_STAMP_PWDATA[27]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[27]\);
    
    \MemorySynchronizer_0/un1_nreset_49\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[6]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_nreset_49_i\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_31\ : CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_25_Z\, B
         => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_24_Z\, 
        C => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_23_Z\, 
        D => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_22_Z\, 
        Y => \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_31_Z\);
    
    \STAMP_0/measurement_dms1_0_sqmuxa_1_1_a3\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \STAMP_0/apb_spi_finished_0_sqmuxa_1\, B => 
        debug_led_net_0, C => \STAMP_0/spi_request_for_Z[1]\, D
         => \STAMP_0/spi_request_for_Z[0]\, Y => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\);
    
    \MemorySynchronizer_0/resynctimercounter[30]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1092\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[30]\);
    
    \STAMP_0/drdy_flank_detected_temp_RNO\ : CFG1
      generic map(INIT => "01")

      port map(A => stamp0_ready_temp_c, Y => 
        \STAMP_0/stamp0_ready_temp_c_i\);
    
    \STAMP_0/spi/clk_toggles_cry[1]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/spi/clk_toggles_Z[1]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/spi/clk_toggles_s_390_FCO\, S
         => \STAMP_0/spi/clk_toggles_s[1]\, Y => OPEN, FCO => 
        \STAMP_0/spi/clk_toggles_cry_Z[1]\, CC => 
        NET_CC_CONFIG610, P => NET_CC_CONFIG608, UB => 
        NET_CC_CONFIG609);
    
    AFLSDF_INV_78 : INV_BA
      port map(A => debug_led_net_0, Y => \AFLSDF_INV_78\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[7]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_7_S\, 
        Y => \MemorySynchronizer_0/N_1545\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_47\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1]\, 
        IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data_0[13]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[13]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[13]\, Y
         => \STAMP_0/N_596\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a0_1\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => \MemorySynchronizer_0/N_2313\, C => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_29_Z\, 
        D => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_a2_0_32_30_Z\, 
        Y => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_0_a0_1_Z\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_45_set_RNI93UF\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_45_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[27]\, C
         => \MemorySynchronizer_0/un1_nreset_38_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[27]\);
    
    \STAMP_0/spi/tx_buffer[9]\ : SLE
      port map(D => \STAMP_0/spi/N_126\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[9]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_221\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10[16]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/ConfigReg_Z[16]\, B => 
        \MemorySynchronizer_0/N_2567\, C => 
        \MemorySynchronizer_0/N_2586\, Y => 
        \MemorySynchronizer_0/N_1228\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_27\ : CFG4
      generic map(INIT => x"1000")

      port map(A => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_25_S\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_24_S\, 
        C => \MemorySynchronizer_0/un6_in_enable_0_a3_23_Z\, D
         => \MemorySynchronizer_0/un6_in_enable_0_a3_13_Z\, Y => 
        \MemorySynchronizer_0/un6_in_enable_0_a3_27_Z\);
    
    \MemorySynchronizer_0/un1_nreset_23\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[10]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_23_i\);
    
    \STAMP_0/drdy_flank_detected_dms2_RNO\ : CFG1
      generic map(INIT => "01")

      port map(A => stamp0_ready_dms2_c, Y => 
        \STAMP_0/stamp0_ready_dms2_c_i\);
    
    \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc0\ : 
        CFG4
      generic map(INIT => x"338C")

      port map(A => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[1]\, B => 
        \MemorySynchronizer_0/enableTimestampGen_Z\, C => 
        \MemorySynchronizer_0/TimeStampGen/un6_enable_3_Z\, D => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[0]\, Y => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc0_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg[26]\ : SLE
      port map(D => \MemorySynchronizer_0/N_2034_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[26]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_249\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[2]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_2\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[16]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[16]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[16]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[16]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[16]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[3]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[3]\);
    
    \MemorySynchronizer_0/un1_nreset_3_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[11]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_3_i\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_218\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_40_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_92\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_40_set_Z\);
    
    \STAMP_0/measurement_dms1[9]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[57]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_36_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_93\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_36_set_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[22]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[1]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[22]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[22]\);
    
    \MemorySynchronizer_0/TimeStampGen/prescaler_5[3]\ : CFG4
      generic map(INIT => x"1230")

      port map(A => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_c2\, B
         => \MemorySynchronizer_0/TimeStampGen/countere\, C => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[3]\, D => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[2]\, Y => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_5_Z[3]\);
    
    \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa_0_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0080")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[3]\, 
        B => ENABLE_MEMORY_LED_c, C => 
        \MemorySynchronizer_0/N_140_2\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[29]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_29\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[29]\, 
        C => \MemorySynchronizer_0/N_1480\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[29]\);
    
    \MemorySynchronizer_0/resettimercounter[9]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[9]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_44_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[9]\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_24\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/N_1084\, B => 
        \MemorySynchronizer_0/N_1081\, C => 
        \MemorySynchronizer_0/N_1068\, D => 
        \MemorySynchronizer_0/N_1065\, Y => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_24_Z\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_37_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_94\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_37_set_Z\);
    
    \adc_start_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \adc_start_obuf/U0/DOUT1\, Y => 
        \adc_start_obuf/U0/DOUT\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_55\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[6]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[6]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[6]\, C => 
        \MemorySynchronizer_0/N_2593\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[6]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[15]\ : SLE
      port map(D => \STAMP_0_data_frame[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[15]\);
    
    AFLSDF_INV_52 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_58_Z\, Y => 
        \AFLSDF_INV_52\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[16]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[16]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[16]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_0_a1_1\ : 
        CFG3
      generic map(INIT => x"08")

      port map(A => \MemorySynchronizer_0/APBState_Z[0]\, B => 
        \sb_sb_0_STAMP_PADDR[3]\, C => \sb_sb_0_STAMP_PADDR[6]\, 
        Y => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_0_a1_1_Z\);
    
    \LED_HEARTBEAT_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => LED_HEARTBEAT, D => 
        \LED_HEARTBEAT_obuf/U0/DOUT\, E => 
        \LED_HEARTBEAT_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[30]\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_0_Z[30]\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[30]\, C => 
        \MemorySynchronizer_0/N_2593\, D => 
        \MemorySynchronizer_0/N_1217\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[30]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_75\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16]\, 
        IPC => OPEN);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[1]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[1]\, B => 
        \sb_sb_0_Memory_PRDATA[1]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1]\);
    
    AFLSDF_INV_15 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_60\, Y => 
        \AFLSDF_INV_15\);
    
    \STAMP_0/spi/count[28]\ : SLE
      port map(D => \STAMP_0/spi/count_lm[28]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_49_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi/count_Z[28]\);
    
    \STAMP_0/spi/un7_count_NE_20\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \STAMP_0/spi/count_Z[3]\, B => 
        \STAMP_0/spi/count_Z[2]\, C => \STAMP_0/spi/count_Z[1]\, 
        D => \STAMP_0/spi/count_Z[0]\, Y => 
        \STAMP_0/spi/un7_count_NE_20_Z\);
    
    \STAMP_0/spi/tx_buffer_RNO[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[14]\, B => 
        \STAMP_0/spi/tx_buffer_Z[13]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_121\);
    
    \MOSI_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => MOSI, D => \MOSI_obuf/U0/DOUT\, E => 
        \MOSI_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[5]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[5]\, B => 
        \sb_sb_0_STAMP_PWDATA[5]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[5]\);
    
    \MemorySynchronizer_0/SynchronizerInterrupt_RNO\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \MemorySynchronizer_0/N_2567\, B => 
        \MemorySynchronizer_0/N_2586\, C => 
        \MemorySynchronizer_0/APBState_Z[1]\, D => 
        \sb_sb_0_STAMP_PWDATA[30]\, Y => 
        \MemorySynchronizer_0/SynchronizerInterrupt_0_sqmuxa_i\);
    
    \STAMP_0/config[4]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[4]\);
    
    \MemorySynchronizer_0/un1_nreset_10_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_37_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_10_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_10_rs_Z\);
    
    \STAMP_0/spi/count_cry[12]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[12]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[11]\, S => 
        \STAMP_0/spi/count_s[12]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[12]\, CC => NET_CC_CONFIG961, P
         => NET_CC_CONFIG959, UB => NET_CC_CONFIG960);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[19]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[19]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[19]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[13]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[19]\);
    
    AFLSDF_INV_103 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_103\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_29_RNI3CT6A\ : 
        CFG4
      generic map(INIT => x"070F")

      port map(A => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_28_Z\, 
        B => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_29_Z\, 
        C => STAMP_0_new_avail, D => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[15]\, Y
         => \MemorySynchronizer_0/N_140_i_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[12]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[12]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[12]\, C => 
        \MemorySynchronizer_0/N_2598\, D => 
        \MemorySynchronizer_0/N_2576\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[12]\);
    
    \STAMP_0/spi/count_lm_0[4]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[4]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[4]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[23]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_23_S\, 
        Y => \MemorySynchronizer_0/N_1505\);
    
    \MemorySynchronizer_0/resynctimercounter[15]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1107\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[15]\);
    
    \MemorySynchronizer_0/un1_nreset_7_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_35_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_7_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_7_rs_Z\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[2]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[2]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_88\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[4]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_26_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_51\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_26_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_26_rs_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[20]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[20]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[19]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[20]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[20]\, CC
         => NET_CC_CONFIG66, P => NET_CC_CONFIG64, UB => 
        NET_CC_CONFIG65);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[21]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[21]\, 
        B => \MemorySynchronizer_0/SynchStatusReg_Z[23]\, C => 
        \MemorySynchronizer_0/N_1182\, D => 
        \MemorySynchronizer_0/N_2580\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[21]\);
    
    \STAMP_0/spi/tx_buffer[13]\ : SLE
      port map(D => \STAMP_0/spi/N_122\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[13]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_28\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[28]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_27_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_28_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_28_Z\, CC
         => NET_CC_CONFIG809, P => NET_CC_CONFIG807, UB => 
        NET_CC_CONFIG808);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3[6]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => \MemorySynchronizer_0/N_2597\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[6]\, C => 
        \MemorySynchronizer_0/TimeStampReg_Z[6]\, D => 
        \MemorySynchronizer_0/N_1254\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[6]\);
    
    
        \MemorySynchronizer_0/copy_and_mark_data.un151_in_enablelto30_13\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/temp_1[5]\, B => 
        \MemorySynchronizer_0/temp_1[6]\, C => 
        \MemorySynchronizer_0/temp_1[7]\, D => 
        \MemorySynchronizer_0/temp_1[8]\, Y => 
        \MemorySynchronizer_0/un151_in_enablelto30_13\);
    
    \MemorySynchronizer_0/PRDATA[30]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21[30]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[30]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[15]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[15]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[15]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[0]\ : SLE
      port map(D => \STAMP_0_data_frame[32]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[0]\);
    
    \STAMP_0/measurement_temp[0]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[16]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_33\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_5\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[5]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_4_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_i_A[5]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_5_Z\, 
        CC => NET_CC_CONFIG119, P => NET_CC_CONFIG117, UB => 
        NET_CC_CONFIG118);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_0\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_1\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => ADLIB_GND0, S => OPEN, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_0_Z\, 
        CC => NET_CC_CONFIG1023, P => NET_CC_CONFIG1021, UB => 
        NET_CC_CONFIG1022);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_1_CC_1\ : CC_CONFIG
      port map(CI => CI_TO_CO535, CO => OPEN, P(0) => 
        NET_CC_CONFIG560, P(1) => NET_CC_CONFIG563, P(2) => 
        NET_CC_CONFIG566, P(3) => NET_CC_CONFIG569, P(4) => 
        NET_CC_CONFIG572, P(5) => NET_CC_CONFIG575, P(6) => 
        NET_CC_CONFIG578, P(7) => NET_CC_CONFIG581, P(8) => 
        NET_CC_CONFIG584, P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, 
        P(11) => ADLIB_VCC1, UB(0) => NET_CC_CONFIG561, UB(1) => 
        NET_CC_CONFIG564, UB(2) => NET_CC_CONFIG567, UB(3) => 
        NET_CC_CONFIG570, UB(4) => NET_CC_CONFIG573, UB(5) => 
        NET_CC_CONFIG576, UB(6) => NET_CC_CONFIG579, UB(7) => 
        NET_CC_CONFIG582, UB(8) => NET_CC_CONFIG585, UB(9) => 
        ADLIB_VCC1, UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, 
        CC(0) => NET_CC_CONFIG562, CC(1) => NET_CC_CONFIG565, 
        CC(2) => NET_CC_CONFIG568, CC(3) => NET_CC_CONFIG571, 
        CC(4) => NET_CC_CONFIG574, CC(5) => NET_CC_CONFIG577, 
        CC(6) => NET_CC_CONFIG580, CC(7) => NET_CC_CONFIG583, 
        CC(8) => NET_CC_CONFIG586, CC(9) => nc359, CC(10) => 
        nc204, CC(11) => nc173);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4[7]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[7]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[7]\, C => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[7]\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_20\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_21\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_19_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[21]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_20_Z\, CC
         => NET_CC_CONFIG1083, P => NET_CC_CONFIG1081, UB => 
        NET_CC_CONFIG1082);
    
    \MemorySynchronizer_0/TimeStampReg[30]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[30]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[30]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_192\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20]\);
    
    \STAMP_0/un1_spi_rx_data_1[7]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[39]\, B => 
        \STAMP_0/dummy_Z[7]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_624\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[23]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[23]\, B => 
        \sb_sb_0_Memory_PRDATA[23]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[23]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_251\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3]\, 
        IPC => OPEN);
    
    \STAMP_0/un52_paddr_5\ : CFG2
      generic map(INIT => x"1")

      port map(A => \sb_sb_0_STAMP_PADDR[3]\, B => 
        \sb_sb_0_STAMP_PADDR[2]\, Y => \STAMP_0/un52_paddr_5_Z\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[18]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[18]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_44\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net\, IPC
         => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter[12]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[12]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_54_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[12]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[6]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[6]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[5]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[6]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[6]\, CC
         => NET_CC_CONFIG24, P => NET_CC_CONFIG22, UB => 
        NET_CC_CONFIG23);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[13]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[13]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[19]\, Y
         => \MemorySynchronizer_0/N_1078\);
    
    \STAMP_0/delay_counter_RNIKM2J[10]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \STAMP_0/delay_counter_Z[11]\, B => 
        \STAMP_0/delay_counter_Z[10]\, C => 
        \STAMP_0/delay_counter_Z[9]\, D => 
        \STAMP_0/delay_counter_Z[8]\, Y => 
        \STAMP_0/N_517_i_0_a2_16\);
    
    \STAMP_0/config[21]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[21]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[21]\);
    
    \MemorySynchronizer_0/un1_nreset_13_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_40_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_13_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_13_rs_Z\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_26\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_27\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_25_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[27]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_26_Z\, CC
         => NET_CC_CONFIG1101, P => NET_CC_CONFIG1099, UB => 
        NET_CC_CONFIG1100);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_12\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[12]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_11_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[20]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_12_Z\, CC
         => NET_CC_CONFIG333, P => NET_CC_CONFIG331, UB => 
        NET_CC_CONFIG332);
    
    \SCLK_obuf/U0/U_IOOUTFF\ : IOOUTFF_BYPASS
      port map(A => \SCLK_obuf/U0/DOUT1\, Y => 
        \SCLK_obuf/U0/DOUT\);
    
    \STAMP_0/un1_async_prescaler_countlto11\ : CFG4
      generic map(INIT => x"0F4F")

      port map(A => \STAMP_0/async_prescaler_count_Z[9]\, B => 
        \STAMP_0/un1_async_prescaler_countlt10\, C => 
        \STAMP_0/async_prescaler_count_Z[11]\, D => 
        \STAMP_0/async_prescaler_count_Z[10]\, Y => 
        \STAMP_0/un1_async_prescaler_count\);
    
    \STAMP_0/spi_tx_data[4]\ : SLE
      port map(D => \STAMP_0/N_294_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[4]\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_16\ : 
        CFG4
      generic map(INIT => x"0004")

      port map(A => \MemorySynchronizer_0/un104_in_enable_axb_31\, 
        B => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_Y\, C
         => \MemorySynchronizer_0/un120_in_enable_i_A[1]\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[30]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_16_Z\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[14]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[14]\);
    
    \MemorySynchronizer_0/TimeStampReg[24]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[24]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[24]\);
    
    \MemorySynchronizer_0/MemorySyncState_RNICHGB[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => ENABLE_MEMORY_LED_c, B => 
        \MemorySynchronizer_0/MemorySyncState_Z[0]\, Y => 
        \MemorySynchronizer_0/N_2028_i\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv[17]\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_17\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[17]\, 
        C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[14]\, D
         => \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, 
        Y => \MemorySynchronizer_0/waitingtimercounter_10[17]\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_5\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[5]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[5]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_4\, S => 
        \MemorySynchronizer_0/temp_1[5]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_5\, CC => 
        NET_CC_CONFIG214, P => NET_CC_CONFIG212, UB => 
        NET_CC_CONFIG213);
    
    \MemorySynchronizer_0/un1_nreset_33_rs_RNIF3FB\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_2537_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[1]\, C => 
        \MemorySynchronizer_0/un1_nreset_33_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[1]\);
    
    AFLSDF_INV_94 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_37_Z\, Y => 
        \AFLSDF_INV_94\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_51\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[2]\, B => NN_1, 
        Y => \MemorySynchronizer_0/un1_ResetTimerValueReg_51_Z\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_26\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[26]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_25_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_26_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_26_Z\, 
        CC => NET_CC_CONFIG705, P => NET_CC_CONFIG703, UB => 
        NET_CC_CONFIG704);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_15\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[15]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[15]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_14\, S => 
        \MemorySynchronizer_0/temp_1[15]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_15\, CC => 
        NET_CC_CONFIG244, P => NET_CC_CONFIG242, UB => 
        NET_CC_CONFIG243);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[27]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[27]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[26]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[27]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[27]\, CC
         => NET_CC_CONFIG87, P => NET_CC_CONFIG85, UB => 
        NET_CC_CONFIG86);
    
    \STAMP_0/PRDATA[10]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[10]\);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_23\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/N_1087\, B => 
        \MemorySynchronizer_0/N_1083\, C => 
        \MemorySynchronizer_0/N_1070\, D => 
        \MemorySynchronizer_0/N_1067\, Y => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_23_Z\);
    
    \MemorySynchronizer_0/un1_nreset_61_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_33_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_61_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_61_rs_Z\);
    
    \STAMP_0/un5_async_prescaler_count_cry_10\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[10]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_9_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_10_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_10_Z\, CC
         => NET_CC_CONFIG510, P => NET_CC_CONFIG508, UB => 
        NET_CC_CONFIG509);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO[24]\ : CFG4
      generic map(INIT => x"0F0B")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[24]\, 
        B => \MemorySynchronizer_0/MemorySyncState_Z[3]\, C => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_0_a2_0_0_Z[22]\, 
        D => \MemorySynchronizer_0/N_2321\, Y => 
        \MemorySynchronizer_0/N_215_i\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_14\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[14]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_13_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[18]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_14_Z\, CC
         => NET_CC_CONFIG339, P => NET_CC_CONFIG337, UB => 
        NET_CC_CONFIG338);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7[21]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[21]\, B => 
        \MemorySynchronizer_0/un104_in_enable_21\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[21]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[25]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[25]\);
    
    \STAMP_0/spi/un7_count_NE_21\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \STAMP_0/spi/count_Z[31]\, B => 
        \STAMP_0/spi/count_Z[30]\, C => \STAMP_0/spi/count_Z[29]\, 
        D => \STAMP_0/spi/count_Z[28]\, Y => 
        \STAMP_0/spi/un7_count_NE_21_Z\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS[2]\ : CFG4
      generic map(INIT => x"20A0")

      port map(A => \sb_sb_0/STAMP_PADDRS[14]\, B => 
        \sb_sb_0/STAMP_PADDRS[13]\, C => 
        \sb_sb_0/CoreAPB3_0/iPSELS_raw_1_0_Z[0]\, D => 
        \sb_sb_0/STAMP_PADDRS[12]\, Y => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS_Z[2]\);
    
    \MemorySynchronizer_0/un1_nreset_30_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_58_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_30_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_30_rs_Z\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[16]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[16]\);
    
    \STAMP_0/un1_async_prescaler_countlto8\ : CFG4
      generic map(INIT => x"DFFF")

      port map(A => \STAMP_0/async_prescaler_count_Z[6]\, B => 
        \STAMP_0/un1_async_prescaler_countlt8\, C => 
        \STAMP_0/async_prescaler_count_Z[8]\, D => 
        \STAMP_0/async_prescaler_count_Z[7]\, Y => 
        \STAMP_0/un1_async_prescaler_countlt10\);
    
    \STAMP_0/spi/tx_buffer[3]\ : SLE
      port map(D => \STAMP_0/spi/N_136\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[3]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[17]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[17]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[29]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_29_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[3]\);
    
    \STAMP_0/un1_spi_rx_data_0[10]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[10]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[10]\, Y
         => \STAMP_0/N_593\);
    
    \MemorySynchronizer_0/waitingtimercounter[4]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[4]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_4_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[4]\);
    
    \sb_sb_0/CoreAPB3_0/iPSELS_raw[6]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \sb_sb_0/STAMP_PADDRS[14]\, B => 
        \sb_sb_0/STAMP_PADDRS[13]\, C => 
        \sb_sb_0/CoreAPB3_0/iPSELS_raw_1_0_Z[0]\, D => 
        \sb_sb_0/STAMP_PADDRS[12]\, Y => sb_sb_0_Memory_PSELx);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_34_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_95\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_34_set_Z\);
    
    \MemorySynchronizer_0/ConfigReg_RNO[30]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \sb_sb_0_STAMP_PWDATA[30]\, B => 
        \MemorySynchronizer_0/APBState_Z[1]\, Y => 
        \MemorySynchronizer_0/N_2306_i\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_s[31]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[31]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[30]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s_Z[31]\, 
        Y => OPEN, FCO => OPEN, CC => NET_CC_CONFIG99, P => 
        NET_CC_CONFIG97, UB => NET_CC_CONFIG98);
    
    \STAMP_0/delay_counter_cry[0]_CC_2\ : CC_CONFIG
      port map(CI => CI_TO_CO392, CO => OPEN, P(0) => 
        NET_CC_CONFIG465, P(1) => NET_CC_CONFIG468, P(2) => 
        NET_CC_CONFIG471, P(3) => NET_CC_CONFIG474, P(4) => 
        ADLIB_VCC1, P(5) => ADLIB_VCC1, P(6) => ADLIB_VCC1, P(7)
         => ADLIB_VCC1, P(8) => ADLIB_VCC1, P(9) => ADLIB_VCC1, 
        P(10) => ADLIB_VCC1, P(11) => ADLIB_VCC1, UB(0) => 
        NET_CC_CONFIG466, UB(1) => NET_CC_CONFIG469, UB(2) => 
        NET_CC_CONFIG472, UB(3) => NET_CC_CONFIG475, UB(4) => 
        ADLIB_VCC1, UB(5) => ADLIB_VCC1, UB(6) => ADLIB_VCC1, 
        UB(7) => ADLIB_VCC1, UB(8) => ADLIB_VCC1, UB(9) => 
        ADLIB_VCC1, UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, 
        CC(0) => NET_CC_CONFIG467, CC(1) => NET_CC_CONFIG470, 
        CC(2) => NET_CC_CONFIG473, CC(3) => NET_CC_CONFIG476, 
        CC(4) => nc278, CC(5) => nc169, CC(6) => nc423, CC(7) => 
        nc78, CC(8) => nc263, CC(9) => nc335, CC(10) => nc24, 
        CC(11) => nc409);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_173\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un104_in_enable_cry_0_CC_1\ : CC_CONFIG
      port map(CI => CI_TO_CO819, CO => CI_TO_CO820, P(0) => 
        NET_CC_CONFIG857, P(1) => NET_CC_CONFIG860, P(2) => 
        NET_CC_CONFIG863, P(3) => NET_CC_CONFIG866, P(4) => 
        NET_CC_CONFIG869, P(5) => NET_CC_CONFIG872, P(6) => 
        NET_CC_CONFIG875, P(7) => NET_CC_CONFIG878, P(8) => 
        NET_CC_CONFIG881, P(9) => NET_CC_CONFIG884, P(10) => 
        NET_CC_CONFIG887, P(11) => NET_CC_CONFIG890, UB(0) => 
        NET_CC_CONFIG858, UB(1) => NET_CC_CONFIG861, UB(2) => 
        NET_CC_CONFIG864, UB(3) => NET_CC_CONFIG867, UB(4) => 
        NET_CC_CONFIG870, UB(5) => NET_CC_CONFIG873, UB(6) => 
        NET_CC_CONFIG876, UB(7) => NET_CC_CONFIG879, UB(8) => 
        NET_CC_CONFIG882, UB(9) => NET_CC_CONFIG885, UB(10) => 
        NET_CC_CONFIG888, UB(11) => NET_CC_CONFIG891, CC(0) => 
        NET_CC_CONFIG859, CC(1) => NET_CC_CONFIG862, CC(2) => 
        NET_CC_CONFIG865, CC(3) => NET_CC_CONFIG868, CC(4) => 
        NET_CC_CONFIG871, CC(5) => NET_CC_CONFIG874, CC(6) => 
        NET_CC_CONFIG877, CC(7) => NET_CC_CONFIG880, CC(8) => 
        NET_CC_CONFIG883, CC(9) => NET_CC_CONFIG886, CC(10) => 
        NET_CC_CONFIG889, CC(11) => NET_CC_CONFIG892);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[10]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_10_S\, 
        Y => \MemorySynchronizer_0/N_2434\);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO_3[5]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \MemorySynchronizer_0/numberofnewavails_Z[2]\, 
        B => \MemorySynchronizer_0/m3_e_0_0\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/N_140_2\, Y => 
        \MemorySynchronizer_0/g3\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[24]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[24]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[24]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[8]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[24]\);
    
    \STAMP_0/spi/count_lm_0[22]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[22]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[22]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[19]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[3]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[19]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[19]\);
    
    \MemorySynchronizer_0/TimeStampReg[14]\ : SLE
      port map(D => \MemorySynchronizer_0/TimeStampValue[14]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/N_2304_i\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampReg_Z[14]\);
    
    \MISO_ibuf/U0/U_IOIN\ : IOIN_IB
      port map(YIN => \MISO_ibuf/U0/YIN\, E => ADLIB_GND0, Y => 
        MISO_c);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[8]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[8]\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[7]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[8]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[8]\, CC
         => NET_CC_CONFIG30, P => NET_CC_CONFIG28, UB => 
        NET_CC_CONFIG29);
    
    \STAMP_0/spi/assert_data_RNI4NTB2\ : CFG4
      generic map(INIT => x"44C4")

      port map(A => \STAMP_0/spi/state_Z[0]\, B => 
        \STAMP_0/spi/N_37_i\, C => \STAMP_0/spi/assert_data_Z\, D
         => \STAMP_0/spi/clk_toggles_Z[5]\, Y => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[6]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_6\);
    
    \STAMP_0/spi/tx_buffer_RNO[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[2]\, B => 
        \STAMP_0/spi/tx_buffer_Z[1]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_138\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_a2[10]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \sb_sb_0_STAMP_PADDR[6]\, B => 
        \MemorySynchronizer_0/N_2317\, C => 
        \MemorySynchronizer_0/N_271\, Y => 
        \MemorySynchronizer_0/N_1179\);
    
    \AND2_0_RNIKOS1/U0_RGB1_RGB0\ : RGB_NG
      port map(An => \AND2_0_RNIKOS1/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => OPEN, YR => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB0_rgbr_net_1\);
    
    \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1_0_a2_RNIP7FF\ : 
        CFG2
      generic map(INIT => x"B")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, B => 
        \MemorySynchronizer_0/N_140_1_i\, Y => 
        \MemorySynchronizer_0/N_6\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0_0_0_1[4]\ : CFG4
      generic map(INIT => x"2FAF")

      port map(A => \MemorySynchronizer_0/N_2330\, B => 
        \MemorySynchronizer_0/N_2313\, C => 
        \MemorySynchronizer_0/MemorySyncState_Z[3]\, D => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/MemorySyncState_ns_0_0_0_1_Z[4]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[10]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_10\);
    
    \MemorySynchronizer_0/SynchStatusReg_152_m1_0_0_a2[30]\ : 
        CFG4
      generic map(INIT => x"A0E0")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[2]\, 
        B => \MemorySynchronizer_0/MemorySyncState_Z[0]\, C => 
        ENABLE_MEMORY_LED_c, D => 
        \MemorySynchronizer_0/MemorySyncState_Z[1]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_152_ss0_i_0\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_17\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[17]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[17]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_16\, S => 
        \MemorySynchronizer_0/temp_1[17]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_17\, CC => 
        NET_CC_CONFIG250, P => NET_CC_CONFIG248, UB => 
        NET_CC_CONFIG249);
    
    \MemorySynchronizer_0/SynchStatusReg2[20]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[20]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN
         => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_5_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[20]\);
    
    \STAMP_0/config[29]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[29]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[29]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_53_set_RNI0JNK\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_53_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[13]\, C
         => \MemorySynchronizer_0/un1_nreset_53_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[13]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[26]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[26]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[25]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[26]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[26]\, CC
         => NET_CC_CONFIG84, P => NET_CC_CONFIG82, UB => 
        NET_CC_CONFIG83);
    
    \STAMP_0/spi_dms1_cs_14_iv_i\ : CFG3
      generic map(INIT => x"13")

      port map(A => \STAMP_0/component_state_Z[3]\, B => 
        \STAMP_0/spi_dms1_cs_0_sqmuxa_3\, C => 
        \sb_sb_0_STAMP_PADDR[4]\, Y => 
        \STAMP_0/spi_dms1_cs_14_iv_i_Z\);
    
    \STAMP_0/delay_counter_lm_0[7]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[7]\, Y => 
        \STAMP_0/delay_counter_lm[7]\);
    
    \MemorySynchronizer_0/ConfigReg[25]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[25]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[25]\);
    
    \MemorySynchronizer_0/un1_nreset_33_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_52_i_i_a2_Z\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_33_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_33_rs_Z\);
    
    \STAMP_0/measurement_dms1[7]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[7]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms1_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[55]\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_45_RNIRI17A\ : CFG4
      generic map(INIT => x"0100")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[15]\, B
         => STAMP_0_new_avail, C => \MemorySynchronizer_0/N_6\, D
         => \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, 
        Y => 
        \MemorySynchronizer_0/un112_in_enable_0_I_45_RNIRI17A_Z\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51\ : CFG3
      generic map(INIT => x"08")

      port map(A => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS_Z[2]\, B => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS[1]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PSELSBUS[0]\, Y => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\);
    
    \nCS1_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => nCS1, D => \nCS1_obuf/U0/DOUT\, E => 
        \nCS1_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/un1_nreset_6_rs_RNIDJIR\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_36_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[30]\, C => 
        \MemorySynchronizer_0/un1_nreset_6_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[30]\);
    
    \STAMP_0/un1_spi_rx_data_2[16]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_599\, B => \STAMP_0/N_633\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_666\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[12]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[12]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampValue[12]\);
    
    \MemorySynchronizer_0/un1_nreset_58_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_58_i_i_a2_Z\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_58_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_58_rs_Z\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[7]\ : SLE
      port map(D => \STAMP_0_data_frame[39]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[7]\);
    
    \stamp0_spi_mosi_obuft/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => mosi_1, E => mosi_cl, DOUT => 
        \stamp0_spi_mosi_obuft/U0/DOUT1\, EOUT => 
        \stamp0_spi_mosi_obuft/U0/EOUT1\);
    
    \MemorySynchronizer_0/SynchStatusReg[13]\ : SLE
      port map(D => \MemorySynchronizer_0/SynchStatusReg_168[11]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, 
        EN => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[13]\);
    
    AFLSDF_INV_106 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_44_Z\, Y => 
        \AFLSDF_INV_106\);
    
    AFLSDF_INV_11 : INV_BA
      port map(A => \MemorySynchronizer_0/N_1978_i\, Y => 
        \AFLSDF_INV_11\);
    
    \STAMP_0/spi/tx_buffer_RNO[6]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \STAMP_0/spi_tx_data_Z[6]\, B => 
        \STAMP_0/spi/tx_buffer_Z[5]\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/N_130\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_97\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/COLF_net\, IPB
         => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[3]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_3\);
    
    \STAMP_0/un1_spi_rx_data_2[25]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_608\, B => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, C => \STAMP_0/N_642\, Y
         => \STAMP_0/N_675\);
    
    \STAMP_0/delay_counter_lm_0[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0/N_216_i\, B => 
        \STAMP_0/component_state_RNIFR114_Z[0]\, C => 
        \STAMP_0/delay_counter_s[3]\, Y => 
        \STAMP_0/delay_counter_lm[3]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_19\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[24]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[31]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31]\, 
        IPC => OPEN);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_29\ : 
        CFG4
      generic map(INIT => x"8000")

      port map(A => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_20_Z\, 
        B => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_21_Z\, 
        C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_22_Z\, 
        D => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_23_Z\, 
        Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_29_Z\);
    
    
        \MemorySynchronizer_0/SynchStatusReg_2_sqmuxa_1_0_a2_0_a2_RNIQI741\ : 
        CFG4
      generic map(INIT => x"0054")

      port map(A => STAMP_0_new_avail, B => 
        \MemorySynchronizer_0/N_2028_i\, C => 
        \MemorySynchronizer_0/SynchStatusReg_2_sqmuxa_1\, D => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, Y => 
        \MemorySynchronizer_0/g1\);
    
    \MemorySynchronizer_0/un1_nreset_5_rs_RNIV9221\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_36_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[5]\, C
         => \MemorySynchronizer_0/un1_nreset_5_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[5]\);
    
    \STAMP_0/delay_counter[23]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[23]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[23]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_107\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net\, IPC
         => OPEN);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[11]\ : CFG4
      generic map(INIT => x"0ACE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[11]\, D => 
        \MemorySynchronizer_0/TimeStampReg_Z[11]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[11]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[15]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[15]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[15]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[15]\);
    
    \MMUART_0_TXD_M2F_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => MMUART_0_TXD_M2F_c, E => ADLIB_VCC1, DOUT => 
        \MMUART_0_TXD_M2F_obuf/U0/DOUT1\, EOUT => 
        \MMUART_0_TXD_M2F_obuf/U0/EOUT1\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1[1]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \MemorySynchronizer_0/N_2326\, B => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_1_a2_0_Z[1]\, 
        C => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_0_0_0[4]\, 
        D => \MemorySynchronizer_0/N_2510\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168[1]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[12]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_12_S\, 
        Y => \MemorySynchronizer_0/N_1521\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[11]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_68\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[11]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[11]\, 
        D => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[11]\);
    
    \STAMP_0/spi/count_lm_0[30]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s[30]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[30]\);
    
    \STAMP_0/spi/count_lm_0[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[7]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[7]\);
    
    \sb_sb_0/CCC_0/GL1_INST/U0_RGB1\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL1_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => OPEN, YR => 
        \sb_sb_0/CCC_0/GL1_INST/U0_RGB1_YR\);
    
    \STAMP_0/spi/rx_buffer[4]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[3]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[4]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter[2]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/counter_s[2]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/TimeStampGen/countere\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB8_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/TimeStampValue[2]\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[10]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[10]\, B => 
        \sb_sb_0_Memory_PRDATA[10]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10]\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_17\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/GPD3_ARST_N_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PADDR_net[7]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_33_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_96\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_33_set_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv[22]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, B => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[22]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[22]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_m[10]\, Y
         => \MemorySynchronizer_0/resettimercounter_9[22]\);
    
    \STAMP_0/PRDATA[6]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[6]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_50_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_97\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_50_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_143\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter[13]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[13]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_21_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[13]\);
    
    AFLSDF_INV_45 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_58_i_i_a2_Z\, 
        Y => \AFLSDF_INV_45\);
    
    \STAMP_0/spi/tx_buffer_RNO[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/spi/state_Z[0]\, B => 
        \STAMP_0/spi_tx_data_Z[0]\, Y => \STAMP_0/spi/N_333\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[18]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[18]\, B => 
        \sb_sb_0_Memory_PRDATA[18]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[18]\);
    
    \STAMP_0/un60_paddr_3_2\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \sb_sb_0_STAMP_PADDR[7]\, B => 
        \sb_sb_0_STAMP_PADDR[2]\, C => \sb_sb_0_STAMP_PADDR[3]\, 
        D => \sb_sb_0_STAMP_PADDR[4]\, Y => 
        \STAMP_0/un60_paddr_3_2_Z\);
    
    \STAMP_0/spi_enable_RNO\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/N_361\, B => 
        \STAMP_0/component_state_Z[3]\, Y => 
        \STAMP_0/spi_enable_RNO_Z\);
    
    \STAMP_0/spi/rx_buffer[12]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[12]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[18]\ : SLE
      port map(D => \STAMP_0_data_frame[18]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[18]\);
    
    \STAMP_0/dummy[16]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_98\, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/dummy_Z[16]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_49_set_RNINFNL\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_49_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[24]\, C => 
        \MemorySynchronizer_0/un1_nreset_9_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[24]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[10]\ : SLE
      port map(D => \STAMP_0_data_frame[42]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[10]\);
    
    \STAMP_0/un1_request_resync_0_sqmuxa_1\ : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \STAMP_0/request_resync_0_sqmuxa\, B => 
        \STAMP_0/dummy_1_sqmuxa_2_Z\, C => 
        \STAMP_0/un52_paddr_5_Z\, D => 
        \STAMP_0/dummy_1_sqmuxa_4_Z\, Y => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\);
    
    \STAMP_0/spi/count_lm_0[15]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \STAMP_0/spi/count_s[15]\, B => 
        \STAMP_0/spi/state_Z[0]\, C => 
        \STAMP_0/spi/un7_count_NE_i\, Y => 
        \STAMP_0/spi/count_lm[15]\);
    
    \MemorySynchronizer_0/ResetTimerValueReg[16]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[16]\);
    
    \STAMP_0/un45_async_state_cry_0_CC_0\ : CC_CONFIG
      port map(CI => ADLIB_GND0, CO => OPEN, P(0) => 
        NET_CC_CONFIG514, P(1) => NET_CC_CONFIG517, P(2) => 
        NET_CC_CONFIG520, P(3) => NET_CC_CONFIG523, P(4) => 
        NET_CC_CONFIG526, P(5) => NET_CC_CONFIG529, P(6) => 
        NET_CC_CONFIG532, P(7) => ADLIB_VCC1, P(8) => ADLIB_VCC1, 
        P(9) => ADLIB_VCC1, P(10) => ADLIB_VCC1, P(11) => 
        ADLIB_VCC1, UB(0) => NET_CC_CONFIG515, UB(1) => 
        NET_CC_CONFIG518, UB(2) => NET_CC_CONFIG521, UB(3) => 
        NET_CC_CONFIG524, UB(4) => NET_CC_CONFIG527, UB(5) => 
        NET_CC_CONFIG530, UB(6) => NET_CC_CONFIG533, UB(7) => 
        ADLIB_VCC1, UB(8) => ADLIB_VCC1, UB(9) => ADLIB_VCC1, 
        UB(10) => ADLIB_VCC1, UB(11) => ADLIB_VCC1, CC(0) => 
        NET_CC_CONFIG516, CC(1) => NET_CC_CONFIG519, CC(2) => 
        NET_CC_CONFIG522, CC(3) => NET_CC_CONFIG525, CC(4) => 
        NET_CC_CONFIG528, CC(5) => NET_CC_CONFIG531, CC(6) => 
        NET_CC_CONFIG534, CC(7) => nc88, CC(8) => nc111, CC(9)
         => nc55, CC(10) => nc10, CC(11) => nc22);
    
    \MemorySynchronizer_0/N_2535_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_99\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/N_2535_set_Z\);
    
    AFLSDF_INV_70 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_70\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_7\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[7]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_6_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[25]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_7_Z\, CC
         => NET_CC_CONFIG318, P => NET_CC_CONFIG316, UB => 
        NET_CC_CONFIG317);
    
    \MemorySynchronizer_0/waitingtimercounter_RNI7RIN[18]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_35_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[18]\, C
         => \MemorySynchronizer_0/un1_nreset_46_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[18]\);
    
    \STAMP_0/un5_async_prescaler_count_s_1_391_CC_0\ : CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => CI_TO_CO477, P(0) => 
        ADLIB_VCC1, P(1) => ADLIB_VCC1, P(2) => ADLIB_VCC1, P(3)
         => ADLIB_VCC1, P(4) => ADLIB_VCC1, P(5) => ADLIB_VCC1, 
        P(6) => ADLIB_VCC1, P(7) => ADLIB_VCC1, P(8) => 
        ADLIB_GND0, P(9) => NET_CC_CONFIG478, P(10) => 
        NET_CC_CONFIG481, P(11) => NET_CC_CONFIG484, UB(0) => 
        ADLIB_VCC1, UB(1) => ADLIB_VCC1, UB(2) => ADLIB_VCC1, 
        UB(3) => ADLIB_VCC1, UB(4) => ADLIB_VCC1, UB(5) => 
        ADLIB_VCC1, UB(6) => ADLIB_VCC1, UB(7) => ADLIB_VCC1, 
        UB(8) => ADLIB_GND0, UB(9) => NET_CC_CONFIG479, UB(10)
         => NET_CC_CONFIG482, UB(11) => NET_CC_CONFIG485, CC(0)
         => nc392, CC(1) => nc210, CC(2) => nc185, CC(3) => nc143, 
        CC(4) => nc433, CC(5) => nc417, CC(6) => nc248, CC(7) => 
        nc389, CC(8) => nc77, CC(9) => NET_CC_CONFIG480, CC(10)
         => NET_CC_CONFIG483, CC(11) => NET_CC_CONFIG486);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0_0[11]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[11]\, B => 
        \sb_sb_0_STAMP_PWDATA[11]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[11]\);
    
    \MemorySynchronizer_0/un94_in_enable_20\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/resettimercounter_Z[4]\, 
        B => \MemorySynchronizer_0/resettimercounter_Z[3]\, C => 
        \MemorySynchronizer_0/resettimercounter_Z[2]\, D => 
        \MemorySynchronizer_0/resettimercounter_Z[1]\, Y => 
        \MemorySynchronizer_0/un94_in_enable_20_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[2]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/TimeStampReg_Z[2]\, D => 
        \MemorySynchronizer_0/ConfigReg_Z[2]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[2]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_223\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19]\, 
        IPC => OPEN);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\);
    
    \STAMP_0/delay_counter_cry[23]\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/delay_counter_Z[23]\, C => ADLIB_GND0, D => 
        ADLIB_GND0, FCI => \STAMP_0/delay_counter_cry_Z[22]\, S
         => \STAMP_0/delay_counter_s[23]\, Y => OPEN, FCO => 
        \STAMP_0/delay_counter_cry_Z[23]\, CC => NET_CC_CONFIG464, 
        P => NET_CC_CONFIG462, UB => NET_CC_CONFIG463);
    
    \STAMP_0/config[17]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[17]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[17]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_286\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_28\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[28]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_27_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_28_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_28_Z\, 
        CC => NET_CC_CONFIG711, P => NET_CC_CONFIG709, UB => 
        NET_CC_CONFIG710);
    
    \STAMP_0/spi/rx_buffer[2]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[2]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_29\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[1]\ : SLE
      port map(D => \STAMP_0_data_frame[33]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[1]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[10]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbl_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[10]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_5\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_179\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_a2_1[14]\ : 
        CFG3
      generic map(INIT => x"40")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/N_140_i\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_14_S\, 
        Y => \MemorySynchronizer_0/N_1529\);
    
    \MemorySynchronizer_0/resettimercounter_RNINACO[9]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \MemorySynchronizer_0/N_2535_set_Z\, B => 
        \MemorySynchronizer_0/resettimercounterrs[9]\, C => 
        \MemorySynchronizer_0/un1_nreset_44_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[9]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_175\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[18]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_18\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[18]\, 
        C => \MemorySynchronizer_0/N_1509\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[18]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_0_iv_0_a2_1[31]\ : 
        CFG3
      generic map(INIT => x"04")

      port map(A => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, B
         => \MemorySynchronizer_0/un104_in_enable_axb_31\, C => 
        \MemorySynchronizer_0/N_140_1_i\, Y => 
        \MemorySynchronizer_0/N_2471\);
    
    \STAMP_0/spi/assert_data\ : SLE
      port map(D => \STAMP_0/spi/assert_data_5\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB13_rgbr_net_1\, EN => 
        debug_led_net_0, ALn => ADLIB_VCC1, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \STAMP_0/spi/assert_data_Z\);
    
    \STAMP_0/dummy[11]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB5_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_100\, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/dummy_Z[11]\);
    
    \MemorySynchronizer_0/SynchStatusReg2[0]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/SynchStatusReg2_79_i_i_a2_fast_Z[0]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, 
        EN => 
        \MemorySynchronizer_0/SynchStatusReg2_0_sqmuxa_6_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_10_RNID80A1_Z[31]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[0]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_7\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12]\, 
        IPC => OPEN);
    
    AFLSDF_INV_104 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_104\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[25]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[25]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[25]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[25]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[25]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[25]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_9[4]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[6]\, B
         => \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_16_0_Z[28]\, 
        C => \MemorySynchronizer_0/N_1182\, Y => 
        \MemorySynchronizer_0/N_1260\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_122\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net\, IPB
         => OPEN, IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_282\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9]\, 
        IPC => OPEN);
    
    \STAMP_0/measurement_temp[9]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[25]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_86\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/RXDF_net[2]\, 
        IPC => OPEN);
    
    \STAMP_0/un1_spi_rx_data_1[11]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[43]\, B => 
        \STAMP_0/dummy_Z[11]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_628\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[29]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[29]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[29]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[29]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[28]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_28_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[4]\);
    
    \MemorySynchronizer_0/TimeStampGen/counter_cry[15]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/TimeStampValue[15]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[14]\, S
         => \MemorySynchronizer_0/TimeStampGen/counter_s[15]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/TimeStampGen/counter_cry_Z[15]\, CC
         => NET_CC_CONFIG51, P => NET_CC_CONFIG49, UB => 
        NET_CC_CONFIG50);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_52_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_101\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_52_set_Z\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_3\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_4\, C => ADLIB_GND0, 
        D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_2_Z\, S => 
        \MemorySynchronizer_0/un120_in_enable_a_4[4]\, Y => OPEN, 
        FCO => \MemorySynchronizer_0/un120_in_enable_a_4_cry_3_Z\, 
        CC => NET_CC_CONFIG1032, P => NET_CC_CONFIG1030, UB => 
        NET_CC_CONFIG1031);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO_0[5]\ : CFG4
      generic map(INIT => x"1300")

      port map(A => \MemorySynchronizer_0/N_140_2\, B => 
        \MemorySynchronizer_0/N_6\, C => 
        \MemorySynchronizer_0/N_2330\, D => 
        \MemorySynchronizer_0/SynchStatusReg_RNO_2_Z[5]\, Y => 
        \MemorySynchronizer_0/N_4\);
    
    \MemorySynchronizer_0/PRDATA[16]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21[16]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[16]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_a2_0\ : 
        CFG2
      generic map(INIT => x"4")

      port map(A => \sb_sb_0_STAMP_PADDR[4]\, B => 
        \sb_sb_0_STAMP_PADDR[2]\, Y => 
        \MemorySynchronizer_0/N_2564\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[23]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[23]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[23]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[23]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[17]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[17]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[17]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[17]\);
    
    \STAMP_0/spi_dms1_cs\ : SLE
      port map(D => \STAMP_0/spi_dms1_cs_14_iv_i_Z\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_component_state_14_i_0_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => stamp0_spi_dms1_cs_c);
    
    \MemorySynchronizer_0/SynchStatusReg_RNO[26]\ : CFG4
      generic map(INIT => x"050D")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_4_0_Z[20]\, 
        B => \MemorySynchronizer_0/N_2321\, C => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\, D => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_o2_1_1_Z[20]\, 
        Y => \MemorySynchronizer_0/N_2034_i\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_15[20]\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[31]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[18]\, C => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[14]\, D => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[12]\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_i_i_a2_33_15_Z[20]\);
    
    \MemorySynchronizer_0/MemorySyncState_RNIGLGB[4]\ : CFG2
      generic map(INIT => x"7")

      port map(A => ENABLE_MEMORY_LED_c, B => 
        \MemorySynchronizer_0/MemorySyncState_Z[4]\, Y => 
        \MemorySynchronizer_0/N_2333\);
    
    \STAMP_0/spi/rx_buffer[0]\ : SLE
      port map(D => stamp0_spi_miso_c, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[0]\);
    
    \stamp0_spi_miso_ibuf/U0/U_IOIN\ : IOIN_IB
      port map(YIN => \stamp0_spi_miso_ibuf/U0/YIN\, E => 
        ADLIB_GND0, Y => stamp0_spi_miso_c);
    
    \STAMP_0/un1_spi_rx_data_2[19]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_602\, B => \STAMP_0/N_636\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_669\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0[13]\ : 
        CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[13]\, B => 
        \sb_sb_0_STAMP_PWDATA[13]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[13]\);
    
    \STAMP_0/un1_spi_rx_data_0[28]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame[28]\, B => 
        \STAMP_0/config_Z[28]\, C => \sb_sb_0_STAMP_PADDR[8]\, Y
         => \STAMP_0/N_611\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_225\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_36_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_102\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_36_set_Z\);
    
    \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_o2_0_1[4]\ : 
        CFG4
      generic map(INIT => x"3320")

      port map(A => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_2_0_Z[4]\, 
        B => STAMP_0_new_avail, C => 
        \MemorySynchronizer_0/N_2310\, D => 
        \MemorySynchronizer_0/N_1512\, Y => 
        \MemorySynchronizer_0/N_2509\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1[0]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/SynchStatusReg2_Z[0]\, 
        B => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[0]\, C => 
        \MemorySynchronizer_0/N_2585\, D => 
        \MemorySynchronizer_0/N_2582\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[0]\);
    
    \STAMP_0/spi_request_for_RNO[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/spi_request_for_2_sqmuxa\, B => 
        \STAMP_0/component_state_Z[3]\, Y => \STAMP_0/N_568_i\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_1_CC_0\ : CC_CONFIG
      port map(CI => ADLIB_VCC1, CO => CI_TO_CO535, P(0) => 
        ADLIB_VCC1, P(1) => ADLIB_VCC1, P(2) => ADLIB_VCC1, P(3)
         => ADLIB_GND0, P(4) => NET_CC_CONFIG536, P(5) => 
        NET_CC_CONFIG539, P(6) => NET_CC_CONFIG542, P(7) => 
        NET_CC_CONFIG545, P(8) => NET_CC_CONFIG548, P(9) => 
        NET_CC_CONFIG551, P(10) => NET_CC_CONFIG554, P(11) => 
        NET_CC_CONFIG557, UB(0) => ADLIB_VCC1, UB(1) => 
        ADLIB_VCC1, UB(2) => ADLIB_VCC1, UB(3) => ADLIB_VCC1, 
        UB(4) => NET_CC_CONFIG537, UB(5) => NET_CC_CONFIG540, 
        UB(6) => NET_CC_CONFIG543, UB(7) => NET_CC_CONFIG546, 
        UB(8) => NET_CC_CONFIG549, UB(9) => NET_CC_CONFIG552, 
        UB(10) => NET_CC_CONFIG555, UB(11) => NET_CC_CONFIG558, 
        CC(0) => nc6, CC(1) => nc109, CC(2) => nc87, CC(3) => 
        nc123, CC(4) => NET_CC_CONFIG538, CC(5) => 
        NET_CC_CONFIG541, CC(6) => NET_CC_CONFIG544, CC(7) => 
        NET_CC_CONFIG547, CC(8) => NET_CC_CONFIG550, CC(9) => 
        NET_CC_CONFIG553, CC(10) => NET_CC_CONFIG556, CC(11) => 
        NET_CC_CONFIG559);
    
    \STAMP_0/spi_tx_data_RNO[14]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \sb_sb_0_STAMP_PWDATA[14]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => \STAMP_0/N_267_i\);
    
    \MemorySynchronizer_0/un120_in_enable_a_4_cry_25\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/un104_in_enable_26\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_24_Z\, S
         => \MemorySynchronizer_0/un120_in_enable_a_4[26]\, Y => 
        OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_a_4_cry_25_Z\, CC
         => NET_CC_CONFIG1098, P => NET_CC_CONFIG1096, UB => 
        NET_CC_CONFIG1097);
    
    \MemorySynchronizer_0/SynchStatusReg[5]\ : SLE
      port map(D => \MemorySynchronizer_0/SynchStatusReg_168[3]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, 
        EN => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_2_i_0_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/SynchStatusReg_Z[5]\);
    
    \STAMP_0/un5_async_prescaler_count_cry_2\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[2]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_1_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_2_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_2_Z\, CC
         => NET_CC_CONFIG486, P => NET_CC_CONFIG484, UB => 
        NET_CC_CONFIG485);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[24]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[24]\, B => 
        \sb_sb_0_Memory_PRDATA[24]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[24]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_67\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_24_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[17]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_24_i\);
    
    \MemorySynchronizer_0/un1_nreset_12_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/N_1980_i\, EN => ADLIB_VCC1, ALn
         => \MemorySynchronizer_0/un1_nreset_12_i\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_12_rs_Z\);
    
    \MemorySynchronizer_0/resettimercounter_RNIOJIK[7]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_46_set_Z\, B
         => \MemorySynchronizer_0/resettimercounterrs[7]\, C => 
        \MemorySynchronizer_0/un1_nreset_48_rs_Z\, Y => 
        \MemorySynchronizer_0/resettimercounter_Z[7]\);
    
    \STAMP_0/measurement_temp[6]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[22]\);
    
    \STAMP_0/PRDATA[18]\ : SLE
      port map(D => \STAMP_0/N_668\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_103\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[18]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_176\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/waitingtimercounter[18]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[18]\, CLK
         => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB10_rgbr_net_1\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_46_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/waitingtimercounterrs[18]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6[31]\ : CFG4
      generic map(INIT => x"FFBA")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[31]\, B => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[31]\, C => 
        \MemorySynchronizer_0/N_2574\, D => 
        \MemorySynchronizer_0/N_1123\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[31]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_253\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_GND0, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13]\, 
        IPC => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1]\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_23\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_28_S\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_29_S\, 
        C => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_30_S\, D
         => \MemorySynchronizer_0/un5_resettimercounter_s_31_S\, 
        Y => \MemorySynchronizer_0/un6_in_enable_0_a3_23_Z\);
    
    AFLSDF_INV_98 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_98\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_274\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_17\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[16]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_17_i\);
    
    \STAMP_0/component_state_ns_0_0_0[1]\ : CFG4
      generic map(INIT => x"0E0A")

      port map(A => \STAMP_0/component_state_Z[4]\, B => 
        \STAMP_0/apb_is_atomic_Z\, C => sb_sb_0_STAMP_PENABLE, D
         => \STAMP_0/component_state_Z[2]\, Y => 
        \STAMP_0/component_state_ns_0_0_0_Z[1]\);
    
    AFLSDF_INV_100 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_100\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[20]\ : SLE
      port map(D => \STAMP_0_data_frame[20]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[20]\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_93\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[17]\, B => 
        \MemorySynchronizer_0/un104_in_enable_16\, C => 
        \MemorySynchronizer_0/un104_in_enable_17\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[16]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[7]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[8]\, CC
         => NET_CC_CONFIG562, P => NET_CC_CONFIG560, UB => 
        NET_CC_CONFIG561);
    
    \MemorySynchronizer_0/un104_in_enable_cry_31_FCINST1\ : 
        FCEND_BUFF_CC
      port map(FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_31_FCNET1\, CO
         => \MemorySynchronizer_0/un104_in_enable_cry_31_Z\, CC
         => NET_CC_CONFIG919, P => NET_CC_CONFIG917, UB => 
        NET_CC_CONFIG918);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[0]\ : SLE
      port map(D => \STAMP_0_data_frame[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB7_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[0]\);
    
    \MemorySynchronizer_0/un112_in_enable_0_I_27\ : ARI1_CC
      generic map(INIT => x"68421")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[15]\, B => 
        \MemorySynchronizer_0/un104_in_enable_14\, C => 
        \MemorySynchronizer_0/un104_in_enable_15\, D => 
        \MemorySynchronizer_0/un120_in_enable_i_A[14]\, FCI => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[6]\, S
         => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[7]\, CC
         => NET_CC_CONFIG559, P => NET_CC_CONFIG557, UB => 
        NET_CC_CONFIG558);
    
    \STAMP_0/un1_spi_rx_data_1[26]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[58]\, B => 
        \STAMP_0/dummy_Z[26]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_643\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \MemorySynchronizer_0/N_1177\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[1]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[1]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[1]\, Y => 
        \MemorySynchronizer_0/PRDATA_21[1]\);
    
    \STAMP_0/PRDATA[20]\ : SLE
      port map(D => \STAMP_0/N_670\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_104\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[20]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_58\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_149\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/ConfigReg[26]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[26]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[26]\);
    
    \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc2\ : 
        CFG2
      generic map(INIT => x"6")

      port map(A => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_c2\, B
         => \MemorySynchronizer_0/TimeStampGen/prescaler_Z[2]\, Y
         => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc2_Z\);
    
    AFLSDF_INV_102 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_36\, Y => 
        \AFLSDF_INV_102\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_145\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/status_dms1_newVal\ : SLE
      port map(D => \STAMP_0/drdy_flank_detected_dms1_0_sqmuxa_1\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, 
        EN => \STAMP_0/un1_drdy_flank_detected_dms1_0_sqmuxa_1_Z\, 
        ALn => \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[15]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[8]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_8\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_21\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[21]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[21]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_20\, S => 
        \MemorySynchronizer_0/temp_1[21]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_21\, CC => 
        NET_CC_CONFIG262, P => NET_CC_CONFIG260, UB => 
        NET_CC_CONFIG261);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_13\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[13]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_12_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_13_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_13_Z\, 
        CC => NET_CC_CONFIG666, P => NET_CC_CONFIG664, UB => 
        NET_CC_CONFIG665);
    
    \STAMP_0/delay_counter[12]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[12]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_152\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_78\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[12]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/un104_in_enable_12\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[14]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[14]\);
    
    \ResetAND_RNIMHJB/U0_RGB1_RGB6\ : RGB_NG
      port map(An => \ResetAND_RNIMHJB/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, YR => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\);
    
    \STAMP_0/un1_spi_rx_data_2[17]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0/N_600\, B => \STAMP_0/N_634\, C => 
        \STAMP_0/un1_spi_rx_data_sn_N_4\, Y => \STAMP_0/N_667\);
    
    \MemorySynchronizer_0/waitingtimercounter[1]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[1]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB9_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_1_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[1]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[29]\ : CFG4
      generic map(INIT => x"0031")

      port map(A => \MemorySynchronizer_0/N_2577\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[29]\, C => 
        \MemorySynchronizer_0/un104_in_enable_29\, D => 
        \MemorySynchronizer_0/N_1403\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[29]\);
    
    \STAMP_0/un1_component_state_9_i_a3\ : CFG3
      generic map(INIT => x"80")

      port map(A => \STAMP_0/un1_component_state_9_i_a3_1_Z\, B
         => \STAMP_0/N_215\, C => \STAMP_0/N_155\, Y => 
        \STAMP_0/N_244\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2_N_2L1_1\ : 
        CFG4
      generic map(INIT => x"EFFF")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[21]\, B => 
        \MemorySynchronizer_0/un120_in_enable_i_A[17]\, C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_21_x_Z\, 
        D => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_20_x_Z\, 
        Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2_N_2L1_1_Z\);
    
    \MemorySynchronizer_0/TimeStampGen/prescaler[0]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc0_Z\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB9_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/TimeStampGen/prescaler_Z[0]\);
    
    AFLSDF_INV_7 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_55\, Y => 
        \AFLSDF_INV_7\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6[10]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[10]\, B => 
        \MemorySynchronizer_0/un104_in_enable_10\, C => 
        \MemorySynchronizer_0/N_2577\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_6_Z[10]\);
    
    \STAMP_0/un1_spi_rx_data_0[15]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame[15]\, B => 
        \sb_sb_0_STAMP_PADDR[8]\, C => \STAMP_0/config_Z[15]\, Y
         => \STAMP_0/N_598\);
    
    \MemorySynchronizer_0/ConfigReg[8]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ConfigReg_0\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/ConfigReg_Z[8]\);
    
    \MemorySynchronizer_0/end_one_counter_0_i_0_o2[0]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => ENABLE_MEMORY_LED_c, B => NN_1, C => 
        \MemorySynchronizer_0/MemorySyncState_Z[1]\, Y => 
        \MemorySynchronizer_0/N_2337\);
    
    \MemorySynchronizer_0/resynctimercounter_1_cry_4\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resynctimercounter_Z[4]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_3_Z\, S
         => \MemorySynchronizer_0/resynctimercounter_1[28]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_4_Z\, CC
         => NET_CC_CONFIG309, P => NET_CC_CONFIG307, UB => 
        NET_CC_CONFIG308);
    
    \STAMP_0/un5_async_prescaler_count_cry_5\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => 
        \STAMP_0/async_prescaler_count_Z[5]\, C => ADLIB_GND0, D
         => ADLIB_GND0, FCI => 
        \STAMP_0/un5_async_prescaler_count_cry_4_Z\, S => 
        \STAMP_0/un5_async_prescaler_count_cry_5_S\, Y => OPEN, 
        FCO => \STAMP_0/un5_async_prescaler_count_cry_5_Z\, CC
         => NET_CC_CONFIG495, P => NET_CC_CONFIG493, UB => 
        NET_CC_CONFIG494);
    
    \STAMP_0/status_async_cycles[5]\ : SLE
      port map(D => \STAMP_0/status_async_cycles_lm[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/status_async_cycles_1_sqmuxa_1_i_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0_data_frame[8]\);
    
    \STAMP_0/config_8_0_a3[31]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \sb_sb_0_STAMP_PWDATA[31]\, B => 
        \STAMP_0/component_state_Z[5]\, Y => 
        \STAMP_0/config_8[31]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_50_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[24]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_50\);
    
    AFLSDF_INV_41 : INV_BA
      port map(A => \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \AFLSDF_INV_41\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0[17]\ : CFG4
      generic map(INIT => x"CC0A")

      port map(A => 
        \MemorySynchronizer_0/waitingtimercounter_Z[17]\, B => 
        \sb_sb_0_STAMP_PWDATA[17]\, C => 
        \MemorySynchronizer_0/N_140_1_i\, D => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, Y
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[17]\);
    
    \STAMP_0/un1_spi_rx_data_0[31]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame[31]\, B => 
        \STAMP_0/config_Z[31]\, C => \sb_sb_0_STAMP_PADDR[8]\, Y
         => \STAMP_0/N_614\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_21\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[21]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_20_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[21]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_21_Z\, 
        CC => NET_CC_CONFIG167, P => NET_CC_CONFIG165, UB => 
        NET_CC_CONFIG166);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_255\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_49_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_56_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_49_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_49_rs_Z\);
    
    \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[8]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \sb_sb_0_STAMP_PRDATA[8]\, B => 
        \sb_sb_0_Memory_PRDATA[8]\, C => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iprdata51_Z\, D => 
        \sb_sb_0/CoreAPB3_0/u_mux_p_to_b3/iPRDATA_0_sqmuxa_Z\, Y
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8]\);
    
    \MemorySynchronizer_0/waitingtimercounter_RNI2V9V[11]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_55_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[11]\, C
         => \MemorySynchronizer_0/un1_nreset_55_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[11]\);
    
    \STAMP_0/spi/count_s[31]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[31]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[30]\, S => 
        \STAMP_0/spi/count_s_Z[31]\, Y => OPEN, FCO => OPEN, CC
         => NET_CC_CONFIG1018, P => NET_CC_CONFIG1016, UB => 
        NET_CC_CONFIG1017);
    
    \MemorySynchronizer_0/resynctimercounter_3_i_0_m2_i_m2[23]\ : 
        CFG3
      generic map(INIT => x"E4")

      port map(A => 
        \MemorySynchronizer_0/resynctimercounter_1_cry_30_Z\, B
         => \MemorySynchronizer_0/resynctimercounter_Z[23]\, C
         => \MemorySynchronizer_0/resynctimercounter_1[9]\, Y => 
        \MemorySynchronizer_0/N_1068\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv[19]\ : CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_19\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_Z[19]\, 
        C => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_m[12]\, D
         => \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, 
        Y => \MemorySynchronizer_0/waitingtimercounter_10[19]\);
    
    \MemorySynchronizer_0/un1_enabletimestampgen2_3_i_a2_0_a2\ : 
        CFG3
      generic map(INIT => x"04")

      port map(A => \MemorySynchronizer_0/MemorySyncState_Z[1]\, 
        B => ENABLE_MEMORY_LED_c, C => 
        \MemorySynchronizer_0/MemorySyncState_Z[0]\, Y => 
        \MemorySynchronizer_0/N_699\);
    
    \MemorySynchronizer_0/waitingtimercounter[0]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/waitingtimercounter_10[0]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_20_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/waitingtimercounterrs[0]\);
    
    \STAMP_0/delay_counter[10]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[10]\);
    
    \MemorySynchronizer_0/un1_nreset_32_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_51_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_32_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_32_rs_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_49\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3]\, 
        IPB => OPEN, IPC => OPEN);
    
    \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11\ : RGB_NG
      port map(An => \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\, ENn
         => ADLIB_GND0, YL => OPEN, YR => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB11_rgbr_net_1\);
    
    \MemorySynchronizer_0/PRDATA[3]\ : SLE
      port map(D => \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[3]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, 
        EN => \MemorySynchronizer_0/APBState_Z[0]\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_Memory_PRDATA[3]\);
    
    \STAMP_0/status_async_cycles_cry[2]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0_data_frame[5]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/status_async_cycles_cry_Z[1]\, S => 
        \STAMP_0/status_async_cycles_s[2]\, Y => OPEN, FCO => 
        \STAMP_0/status_async_cycles_cry_Z[2]\, CC => 
        NET_CC_CONFIG595, P => NET_CC_CONFIG593, UB => 
        NET_CC_CONFIG594);
    
    \MemorySynchronizer_0/WaitingTimerValueReg[9]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \MemorySynchronizer_0/un104_in_enable_9\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_4[31]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \MemorySynchronizer_0/N_2567\, B => 
        \MemorySynchronizer_0/N_271\, C => 
        \MemorySynchronizer_0/ConfigReg_Z[31]\, D => 
        \sb_sb_0_STAMP_PADDR[6]\, Y => 
        \MemorySynchronizer_0/N_1201\);
    
    \STAMP_0/PRDATA[31]\ : SLE
      port map(D => \STAMP_0/N_681\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => \AFLSDF_INV_105\, SD => 
        ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \sb_sb_0_STAMP_PRDATA[31]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_64\ : 
        IP_INTERFACE
      port map(A => ADLIB_GND0, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_281\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_12\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[17]\, B
         => ADLIB_VCC1, C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17]\, 
        IPB => OPEN, IPC => OPEN);
    
    \STAMP_0/spi/count_cry[30]\ : ARI1_CC
      generic map(INIT => x"4AA00")

      port map(A => ADLIB_VCC1, B => \STAMP_0/spi/count_Z[30]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \STAMP_0/spi/count_cry_Z[29]\, S => 
        \STAMP_0/spi/count_s[30]\, Y => OPEN, FCO => 
        \STAMP_0/spi/count_cry_Z[30]\, CC => NET_CC_CONFIG1015, P
         => NET_CC_CONFIG1013, UB => NET_CC_CONFIG1014);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[19]\ : SLE
      port map(D => \STAMP_0_data_frame[19]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[19]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_44_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_106\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_44_set_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_146\ : 
        IP_INTERFACE
      port map(A => RXSM_LO_c, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net\, 
        IPB => OPEN, IPC => OPEN);
    
    \MemorySynchronizer_0/un1_nreset_60_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_60\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_60_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_VCC1, Q => 
        \MemorySynchronizer_0/un1_nreset_60_rs_Z\);
    
    \nCS2_obuf/U0/U_IOTRI\ : IOTRI_OB_EB
      port map(D => nCS2_c, E => ADLIB_VCC1, DOUT => 
        \nCS2_obuf/U0/DOUT1\, EOUT => \nCS2_obuf/U0/EOUT1\);
    
    \MemorySynchronizer_0/resynctimercounter[22]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1100\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[22]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0[13]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_4_Z[13]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_3_Z[13]\, C => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[13]\, D => 
        \MemorySynchronizer_0/N_2574\, Y => 
        \MemorySynchronizer_0/PRDATA_21[13]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_244\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4]\, IPC
         => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_117\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/MemorySyncStatece[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/un6_in_enable_i_0\, B
         => ENABLE_MEMORY_LED_c, C => 
        \MemorySynchronizer_0/MemorySyncState_Z[5]\, Y => 
        \MemorySynchronizer_0/MemorySyncStatece_Z[0]\);
    
    \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_16_0_Z[28]\, B
         => \MemorySynchronizer_0/N_271\, C => 
        \MemorySynchronizer_0/APBState_Z[0]\, D => 
        \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1_0_a2_1_Z\, 
        Y => \MemorySynchronizer_0/SynchStatusReg_1_sqmuxa_1\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_1[1]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \MemorySynchronizer_0/SynchStatusReg_Z[3]\, B
         => \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_16_0_Z[28]\, 
        C => \MemorySynchronizer_0/N_1182\, Y => 
        \MemorySynchronizer_0/N_1172\);
    
    AFLSDF_INV_55 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_44\, Y => 
        \AFLSDF_INV_55\);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_27\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[27]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_26_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_27_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_27_Z\, 
        CC => NET_CC_CONFIG708, P => NET_CC_CONFIG706, UB => 
        NET_CC_CONFIG707);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[10]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_Z[10]\, B => 
        \sb_sb_0_STAMP_PWDATA[10]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D => 
        \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, Y
         => \MemorySynchronizer_0/resettimercounter_9_iv_0_Z[10]\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_38_set_RNI3PRI\ : 
        CFG3
      generic map(INIT => x"EC")

      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_38_set_Z\, 
        B => \MemorySynchronizer_0/waitingtimercounterrs[15]\, C
         => \MemorySynchronizer_0/un1_nreset_51_rs_Z\, Y => 
        \MemorySynchronizer_0/waitingtimercounter_Z[15]\);
    
    \MemorySynchronizer_0/un104_in_enable_cry_26\ : ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/un104_in_enable_26\, B
         => \MemorySynchronizer_0/waitingtimercounter_Z[26]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un104_in_enable_cry_25_Z\, S => 
        OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un104_in_enable_cry_26_Z\, CC => 
        NET_CC_CONFIG901, P => NET_CC_CONFIG899, UB => 
        NET_CC_CONFIG900);
    
    \STAMP_0/config[6]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[6]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[6]\);
    
    \STAMP_0/spi/rx_buffer[10]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/rx_buffer_0_sqmuxa_1\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/spi/rx_buffer_Z[10]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[14]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_14_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[18]\);
    
    \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0[8]\ : 
        CFG4
      generic map(INIT => x"FEFC")

      port map(A => \MemorySynchronizer_0/un104_in_enable_8\, B
         => 
        \MemorySynchronizer_0/waitingtimercounter_10_iv_0_0_0_Z[8]\, 
        C => \MemorySynchronizer_0/N_2430\, D => 
        \MemorySynchronizer_0/waitingtimercounter_3_sqmuxa\, Y
         => \MemorySynchronizer_0/waitingtimercounter_10[8]\);
    
    \MemorySynchronizer_0/resettimercounter[5]\ : SLE
      port map(D => \MemorySynchronizer_0/resettimercounter_9[5]\, 
        CLK => \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, 
        EN => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_50_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => \MemorySynchronizer_0/resettimercounterrs[5]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[24]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[24]\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_Z[24]\, D
         => \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[24]\);
    
    \STAMP_0/delay_counter_RNI6DFR[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \STAMP_0/delay_counter_Z[3]\, B => 
        \STAMP_0/delay_counter_Z[2]\, C => 
        \STAMP_0/delay_counter_Z[1]\, D => 
        \STAMP_0/delay_counter_Z[0]\, Y => 
        \STAMP_0/N_517_i_0_a2_18\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_21\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[21]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_20_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_21_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_21_Z\, CC
         => NET_CC_CONFIG788, P => NET_CC_CONFIG786, UB => 
        NET_CC_CONFIG787);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2[31]\ : CFG4
      generic map(INIT => x"7350")

      port map(A => \MemorySynchronizer_0/Stamp1ShadowReg2_Z[31]\, 
        B => \MemorySynchronizer_0/ResetTimerValueReg_Z[31]\, C
         => \MemorySynchronizer_0/N_2580\, D => 
        \MemorySynchronizer_0/N_2575\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[31]\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_21_x\ : 
        CFG3
      generic map(INIT => x"01")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[18]\, B => 
        \MemorySynchronizer_0/un120_in_enable_i_A[19]\, C => 
        \MemorySynchronizer_0/un120_in_enable_i_A[20]\, Y => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_a2_1_21_x_Z\);
    
    \STAMP_0/spi/un7_count_NE_28\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \STAMP_0/spi/un7_count_NE_19_Z\, B => 
        \STAMP_0/spi/un7_count_NE_18_Z\, C => 
        \STAMP_0/spi/un7_count_NE_17_Z\, D => 
        \STAMP_0/spi/un7_count_NE_16_Z\, Y => 
        \STAMP_0/spi/un7_count_NE_28_Z\);
    
    \STAMP_0/config[24]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[24]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbr_net_1\, EN => 
        \STAMP_0/config_143\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/config_Z[24]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[11]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[11]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[11]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[11]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[11]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[11]\);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_RNO[2]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => 
        \MemorySynchronizer_0/un1_MemorySyncState_11_i\, B => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_2_S\, C
         => \MemorySynchronizer_0/ResetTimerValueReg_1_sqmuxa\, D
         => ENABLE_MEMORY_LED_c, Y => 
        \MemorySynchronizer_0/un5_resettimercounter_m[30]\);
    
    \MemorySynchronizer_0/un6_in_enable_0_a3_21\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_20_S\, B
         => \MemorySynchronizer_0/un5_resettimercounter_cry_21_S\, 
        C => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_22_S\, D
         => \MemorySynchronizer_0/un5_resettimercounter_cry_23_S\, 
        Y => \MemorySynchronizer_0/un6_in_enable_0_a3_21_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[19]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => \MemorySynchronizer_0/TimeStampReg_Z[19]\, B
         => \MemorySynchronizer_0/Stamp1ShadowReg1_Z[19]\, C => 
        \MemorySynchronizer_0/N_2598\, D => 
        \MemorySynchronizer_0/N_2576\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[19]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_49\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[24]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_49_Z\);
    
    \STAMP_0/un1_spi_rx_data[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_653\, C => \STAMP_0/spi_rx_data[3]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[3]\);
    
    \STAMP_0/delay_counter_lm_0[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \STAMP_0/component_state_RNIFR114_Z[0]\, B
         => \STAMP_0/delay_counter_s[5]\, Y => 
        \STAMP_0/delay_counter_lm[5]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_270\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30]\, 
        IPB => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_RREADY_net\, 
        IPC => OPEN);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_11\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/PLL_POWERDOWN_N_net\, IPB
         => \sb_sb_0/CCC_0/CCC_INST/NGMUX3_HOLD_N_net\, IPC => 
        OPEN);
    
    \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_25\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \MemorySynchronizer_0/N_1082\, B => 
        \MemorySynchronizer_0/N_1079\, C => 
        \MemorySynchronizer_0/N_1066\, D => 
        \MemorySynchronizer_0/N_1063\, Y => 
        \MemorySynchronizer_0/un41_in_enable_0_a2_0_a2_25_Z\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_fast[15]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/WaitingTimerValueReg_1_sqmuxa\, ALn
         => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn => 
        ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/WaitingTimerValueReg_fast_Z[15]\);
    
    \STAMP_0/measurement_dms2[12]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[12]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_dms2_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[44]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_121\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net\, IPB
         => OPEN, IPC => OPEN);
    
    \stamp0_spi_temp_cs_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => stamp0_spi_temp_cs, D => 
        \stamp0_spi_temp_cs_obuf/U0/DOUT\, E => 
        \stamp0_spi_temp_cs_obuf/U0/EOUT\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5[0]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \MemorySynchronizer_0/N_2575\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_1_Z[0]\, C => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[0]\, D => 
        \MemorySynchronizer_0/N_1179\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[0]\);
    
    \MemorySynchronizer_0/un4_waitingtimercounter_cry_28\ : 
        ARI1_CC
      generic map(INIT => x"595AA")

      port map(A => \MemorySynchronizer_0/un105_m1_e_0_0\, B => 
        \MemorySynchronizer_0/waitingtimercounter_Z[28]\, C => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_27_Z\, D => 
        \MemorySynchronizer_0/un105_in_enable_i_0_a2_28_Z\, FCI
         => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_27_Z\, 
        S => \MemorySynchronizer_0/un120_in_enable_i_A[28]\, Y
         => OPEN, FCO => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_28_Z\, 
        CC => NET_CC_CONFIG188, P => NET_CC_CONFIG186, UB => 
        NET_CC_CONFIG187);
    
    \STAMP_0/PRDATA[14]\ : SLE
      port map(D => \STAMP_0/un1_spi_rx_data_Z[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_i\, ALn => ADLIB_VCC1, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \sb_sb_0_STAMP_PRDATA[14]\);
    
    \MemorySynchronizer_0/un5_resettimercounter_cry_4\ : ARI1_CC
      generic map(INIT => x"65500")

      port map(A => ADLIB_VCC1, B => 
        \MemorySynchronizer_0/resettimercounter_Z[4]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_3_Z\, S
         => \MemorySynchronizer_0/un5_resettimercounter_cry_4_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un5_resettimercounter_cry_4_Z\, CC
         => NET_CC_CONFIG737, P => NET_CC_CONFIG735, UB => 
        NET_CC_CONFIG736);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[10]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[10]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1081\, Y => 
        \MemorySynchronizer_0/N_1112\);
    
    \STAMP_0/spi/tx_buffer[11]\ : SLE
      port map(D => \STAMP_0/spi/N_124\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB2_rgbr_net_1\, EN => 
        \STAMP_0/spi/un1_reset_n_inv_2_i\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi/tx_buffer_Z[11]\);
    
    \AND2_0_RNIKOS1/U0_RGB1_RGB3\ : RGB_NG
      port map(An => \AND2_0_RNIKOS1/U0_YNn_GSouth\, ENn => 
        ADLIB_GND0, YL => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbl_net_1\, YR => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg2[5]\ : SLE
      port map(D => \STAMP_0_data_frame[5]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_0_sqmuxa_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB4_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_13_RNILNGL_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg2_Z[5]\);
    
    \MemorySynchronizer_0/un1_nreset_37_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[28]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_37_i\);
    
    \sb_sb_0/CCC_0/CCC_INST/IP_INTERFACE_2\ : IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => \sb_sb_0/CCC_0/CCC_INST/PCLK_net\, IPB => 
        \sb_sb_0/CCC_0/CCC_INST/NGMUX0_SEL_net\, IPC => 
        \sb_sb_0/CCC_0/CCC_INST/PWDATA_net[0]\);
    
    \STAMP_0/spi_tx_data[3]\ : SLE
      port map(D => \STAMP_0/N_295_i\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbl_net_1\, EN => 
        \STAMP_0/un1_presetn_inv_2_i_0_Z\, ALn => ADLIB_VCC1, ADn
         => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => \STAMP_0/spi_tx_data_Z[3]\);
    
    \STAMP_0/un1_spi_rx_data_1[29]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[61]\, B => 
        \STAMP_0/dummy_Z[29]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_646\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_22\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_29\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => 
        \MemorySynchronizer_0/un120_in_enable_i_A[29]\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_data_tmp[15]\, C
         => ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_28_Z\, 
        S => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_29_S\, 
        Y => OPEN, FCO => 
        \MemorySynchronizer_0/un1_waitingtimercounter_1_cry_29_Z\, 
        CC => NET_CC_CONFIG714, P => NET_CC_CONFIG712, UB => 
        NET_CC_CONFIG713);
    
    \MemorySynchronizer_0/resynctimercounter_5_i_m2_i_m2[28]\ : 
        CFG3
      generic map(INIT => x"E2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[28]\, B => 
        \MemorySynchronizer_0/N_2315\, C => 
        \MemorySynchronizer_0/N_1063\, Y => 
        \MemorySynchronizer_0/N_1094\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_48_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB6_rgbl_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_107\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_48_set_Z\);
    
    \MemorySynchronizer_0/resettimercounter_9_0_iv_0[31]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => 
        \MemorySynchronizer_0/resettimercounter_0_sqmuxa_1\, B
         => \MemorySynchronizer_0/resettimercounter_1_sqmuxa_1\, 
        C => \MemorySynchronizer_0/resettimercounter_Z[31]\, D
         => \MemorySynchronizer_0/un5_resettimercounter_s_31_S\, 
        Y => \MemorySynchronizer_0/resettimercounter_9[31]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_55_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_108\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_55_set_Z\);
    
    \STAMP_0/un27_paddr\ : CFG4
      generic map(INIT => x"CEFF")

      port map(A => \sb_sb_0_STAMP_PADDR[4]\, B => 
        \STAMP_0/un27_paddr_1_Z\, C => stamp0_ready_dms1_c, D => 
        \sb_sb_0_STAMP_PADDR[7]\, Y => \STAMP_0/un27_paddr_i_0\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[17]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[1]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[17]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[17]\);
    
    \MemorySynchronizer_0/SynchStatusReg2_79_fast[13]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \MemorySynchronizer_0/temp_1[2]\, B => 
        \MemorySynchronizer_0/SynchStatusReg2_Z[13]\, C => 
        STAMP_0_new_avail, Y => 
        \MemorySynchronizer_0/SynchStatusReg2_79_fast_Z[13]\);
    
    \MemorySynchronizer_0/un1_nreset_14_rs\ : SLE
      port map(D => ADLIB_VCC1, CLK => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_41_Z\, EN
         => ADLIB_VCC1, ALn => 
        \MemorySynchronizer_0/un1_nreset_14_i\, ADn => ADLIB_VCC1, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_VCC1, Q
         => \MemorySynchronizer_0/un1_nreset_14_rs_Z\);
    
    \MemorySynchronizer_0/resettimercounter[10]\ : SLE
      port map(D => 
        \MemorySynchronizer_0/resettimercounter_9[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB1_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \MemorySynchronizer_0/un1_nreset_23_i\, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resettimercounterrs[10]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_15\ : 
        IP_INTERFACE
      port map(A => 
        \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[20]\, B
         => \sb_sb_0/sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[27]\, 
        C => ADLIB_VCC1, IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27]\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_266\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0]\, 
        IPC => OPEN);
    
    \STAMP_0/un1_presetn_inv_RNIVNUF1\ : CFG2
      generic map(INIT => x"E")

      port map(A => \STAMP_0/un1_presetn_inv_i\, B => 
        \STAMP_0/un1_presetn_inv_RNIK8BR_Z\, Y => 
        \STAMP_0/un1_presetn_inv_RNIVNUF1_Z\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_i[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[3]\, B => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_2_Z[3]\, C => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_5_Z[3]\, D => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_7_Z[3]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_i_Z[3]\);
    
    \STAMP_0/dummy[30]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[30]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_109\, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/dummy_Z[30]\);
    
    \sb_sb_0/CCC_0/GL0_INST\ : GB_NG
      port map(An => \AFLSDF_INV_110\, ENn => ADLIB_GND0, YNn => 
        \sb_sb_0/CCC_0/GL0_INST/U0_YNn\, YSn => 
        \sb_sb_0/CCC_0/GL0_INST/U0_YNn_GSouth\);
    
    \RXSM_SOE_ibuf/U0/U_IOIN\ : IOIN_IB
      port map(YIN => \RXSM_SOE_ibuf/U0/YIN\, E => ADLIB_GND0, Y
         => RXSM_SOE_c);
    
    AFLSDF_INV_22 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_53\, Y => 
        \AFLSDF_INV_22\);
    
    \STAMP_0/spi/rx_data[8]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[8]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[8]\);
    
    \STAMP_0/delay_counter[15]\ : SLE
      port map(D => \STAMP_0/delay_counter_lm[15]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB4_rgbl_net_1\, EN => 
        \STAMP_0/N_118_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB2_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/delay_counter_Z[15]\);
    
    \stamp0_spi_clock_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => stamp0_spi_clock, D => 
        \stamp0_spi_clock_obuf/U0/DOUT\, E => 
        \stamp0_spi_clock_obuf/U0/EOUT\);
    
    AFLSDF_INV_82 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_56_i_i_a2_Z\, 
        Y => \AFLSDF_INV_82\);
    
    \MemorySynchronizer_0/resynctimercounter[28]\ : SLE
      port map(D => \MemorySynchronizer_0/N_1094\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB8_rgbl_net_1\, EN => 
        \MemorySynchronizer_0/N_699\, ALn => 
        \ResetAND_RNIMHJB/U0_RGB1_RGB6_rgbl_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => 
        \MemorySynchronizer_0/resynctimercounter_Z[28]\);
    
    AFLSDF_INV_109 : INV_BA
      port map(A => \STAMP_0/component_state_Z[5]\, Y => 
        \AFLSDF_INV_109\);
    
    \MemorySynchronizer_0/un1_ResyncTimerValueReg_48_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[3]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResyncTimerValueReg_48\);
    
    \stamp0_spi_mosi_obuft/U0/U_IOENFF\ : IOENFF_BYPASS
      port map(A => \stamp0_spi_mosi_obuft/U0/EOUT1\, Y => 
        \stamp0_spi_mosi_obuft/U0/EOUT\);
    
    \STAMP_0/spi/count_lm_0[31]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \STAMP_0/spi/count_s_Z[31]\, B => 
        \STAMP_0/spi/un7_count_NE_i\, C => 
        \STAMP_0/spi/state_Z[0]\, Y => \STAMP_0/spi/count_lm[31]\);
    
    \MemorySynchronizer_0/un1_nreset_60_0_a2_0_a2\ : CFG2
      generic map(INIT => x"E")

      port map(A => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[6]\, B => 
        NN_1, Y => \MemorySynchronizer_0/un1_nreset_60_i\);
    
    \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc1\ : 
        CFG3
      generic map(INIT => x"6C")

      port map(A => \MemorySynchronizer_0/enableTimestampGen_Z\, 
        B => \MemorySynchronizer_0/TimeStampGen/prescaler_Z[1]\, 
        C => \MemorySynchronizer_0/TimeStampGen/prescaler_Z[0]\, 
        Y => 
        \MemorySynchronizer_0/TimeStampGen/un1_prescaler_axbxc1_Z\);
    
    \STAMP_0/spi/rx_data[14]\ : SLE
      port map(D => \STAMP_0/spi/rx_buffer_Z[14]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB3_rgbr_net_1\, EN => 
        \STAMP_0/spi/N_50_i\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB1_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => 
        ADLIB_GND0, Q => \STAMP_0/spi_rx_data[14]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_59_set\ : SLE
      port map(D => CFG0_GND_INST_NET, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB0_rgbr_net_1\, EN => 
        ADLIB_VCC1, ALn => \AFLSDF_INV_111\, ADn => ADLIB_GND0, 
        SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT => ADLIB_GND0, Q
         => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_59_set_Z\);
    
    \MemorySynchronizer_0/MemorySyncState_ns_0[0]\ : CFG4
      generic map(INIT => x"ABAA")

      port map(A => 
        \MemorySynchronizer_0/MemorySyncState_ns_0_1_Z[0]\, B => 
        STAMP_0_new_avail, C => 
        \MemorySynchronizer_0/un41_in_enable_i_0\, D => 
        \MemorySynchronizer_0/N_1495\, Y => 
        \MemorySynchronizer_0/MemorySyncState_ns[0]\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[6]\ : SLE
      port map(D => \STAMP_0_data_frame[38]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[6]\);
    
    \MemorySynchronizer_0/ResyncTimerValueReg[11]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[11]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/ResyncTimerValueReg_1_sqmuxa_i_i_a2_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB3_rgbr_net_1\, ADn
         => ADLIB_GND0, SLn => ADLIB_VCC1, SD => ADLIB_GND0, LAT
         => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/ResyncTimerValueReg_Z[11]\);
    
    \STAMP_0/dummy[9]\ : SLE
      port map(D => \sb_sb_0_STAMP_PWDATA[9]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/un1_request_resync_0_sqmuxa_1_Z\, ALn => 
        \AND2_0_RNIKOS1/U0_RGB1_RGB3_rgbr_net_1\, ADn => 
        ADLIB_VCC1, SLn => \AFLSDF_INV_112\, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0/dummy_Z[9]\);
    
    \STAMP_0/un85_paddr_3_0_tz\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => \sb_sb_0_STAMP_PADDR[8]\, B => 
        \STAMP_0/un68_paddr_1_0_Z\, C => \sb_sb_0_STAMP_PADDR[9]\, 
        D => \STAMP_0/un60_paddr_3_2_Z\, Y => 
        \STAMP_0/un85_paddr_3_0_tz_Z\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_262\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22]\, 
        IPC => OPEN);
    
    \MemorySynchronizer_0/resettimercounter_9_iv_0[18]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \MemorySynchronizer_0/N_80\, B => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[18]\, C => 
        \MemorySynchronizer_0/resettimercounter_9_iv_0_0_Z[18]\, 
        D => \MemorySynchronizer_0/resettimercounter_2_sqmuxa\, Y
         => \MemorySynchronizer_0/resettimercounter_9[18]\);
    
    \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1[0]\ : CFG4
      generic map(INIT => x"0CAE")

      port map(A => \MemorySynchronizer_0/N_2581\, B => 
        \MemorySynchronizer_0/N_2576\, C => 
        \MemorySynchronizer_0/TimeStampReg_Z[0]\, D => 
        \MemorySynchronizer_0/ConfigReg_Z[0]\, Y => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_0_1_Z[0]\);
    
    \MemorySynchronizer_0/WaitingTimerValueReg_RNIC38O1[0]\ : 
        ARI1_CC
      generic map(INIT => x"62184")

      port map(A => \MemorySynchronizer_0/un120_in_enable_i_A[1]\, 
        B => \MemorySynchronizer_0/un104_in_enable_0\, C => 
        \MemorySynchronizer_0/un104_in_enable_1\, D => 
        \MemorySynchronizer_0/un4_waitingtimercounter_cry_0_Y\, 
        FCI => ADLIB_GND0, S => OPEN, Y => OPEN, FCO => 
        \MemorySynchronizer_0/un120_in_enable_0_data_tmp[0]\, CC
         => NET_CC_CONFIG1117, P => NET_CC_CONFIG1115, UB => 
        NET_CC_CONFIG1116);
    
    \STAMP_0/un1_spi_rx_data[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \STAMP_0/un1_spi_rx_data_sn_N_5\, B => 
        \STAMP_0/N_654\, C => \STAMP_0/spi_rx_data[4]\, Y => 
        \STAMP_0/un1_spi_rx_data_Z[4]\);
    
    \MemorySynchronizer_0/un1_ResetTimerValueReg_34\ : CFG2
      generic map(INIT => x"2")

      port map(A => 
        \MemorySynchronizer_0/ResetTimerValueReg_Z[29]\, B => 
        NN_1, Y => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_34_Z\);
    
    \MemorySynchronizer_0/Stamp1ShadowReg1[4]\ : SLE
      port map(D => \STAMP_0_data_frame[36]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB7_rgbr_net_1\, EN => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_0_sqmuxa_1_i_0_Z\, 
        ALn => \ResetAND_RNIMHJB/U0_RGB1_RGB5_rgbr_net_1\, ADn
         => ADLIB_VCC1, SLn => 
        \MemorySynchronizer_0/PRDATA_21_0_iv_0_a2_14_0_RNINM1S_Z[28]\, 
        SD => ADLIB_GND0, LAT => ADLIB_GND0, Q => 
        \MemorySynchronizer_0/Stamp1ShadowReg1_Z[4]\);
    
    AFLSDF_INV_33 : INV_BA
      port map(A => 
        \MemorySynchronizer_0/un1_ResetTimerValueReg_57_Z\, Y => 
        \AFLSDF_INV_33\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_240\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_GND0, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52]\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0]\, IPC
         => \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F_WVALID_net\);
    
    
        \MemorySynchronizer_0/un1_waitingtimercounter_1_sqmuxa_i_0_2_RNILIDKC\ : 
        CFG4
      generic map(INIT => x"EAEE")

      port map(A => \MemorySynchronizer_0/g1\, B => 
        \MemorySynchronizer_0/un112_in_enable_0_I_45_RNIRI17A_Z\, 
        C => 
        \MemorySynchronizer_0/numberofnewavails_RNIVL541_1_Z[0]\, 
        D => \MemorySynchronizer_0/N_140_2\, Y => 
        \MemorySynchronizer_0/SynchStatusReg_168_0_iv_0_a2_0_0_0[4]\);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_151\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_VCC1, C => ADLIB_VCC1, 
        IPA => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net\, 
        IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net\, 
        IPC => OPEN);
    
    \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_130\ : 
        IP_INTERFACE
      port map(A => ADLIB_VCC1, B => ADLIB_GND0, C => ADLIB_VCC1, 
        IPA => OPEN, IPB => 
        \sb_sb_0/sb_sb_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12]\, 
        IPC => OPEN);
    
    \STAMP_0/measurement_temp[10]\ : SLE
      port map(D => \STAMP_0/spi_rx_data[10]\, CLK => 
        \sb_sb_0/CCC_0/GL0_INST/U0_RGB1_RGB5_rgbr_net_1\, EN => 
        \STAMP_0/measurement_temp_1_sqmuxa\, ALn => ADLIB_VCC1, 
        ADn => ADLIB_VCC1, SLn => ADLIB_VCC1, SD => ADLIB_GND0, 
        LAT => ADLIB_GND0, Q => \STAMP_0_data_frame[26]\);
    
    \STAMP_0/un1_spi_rx_data_sn_m3\ : CFG3
      generic map(INIT => x"5C")

      port map(A => \sb_sb_0_STAMP_PADDR[8]\, B => 
        \sb_sb_0_STAMP_PADDR[7]\, C => \sb_sb_0_STAMP_PADDR[9]\, 
        Y => \STAMP_0/un1_spi_rx_data_sn_N_4\);
    
    \MemorySynchronizer_0/copy_and_mark_data.temp_1_cry_22\ : 
        ARI1_CC
      generic map(INIT => x"5AA55")

      port map(A => \MemorySynchronizer_0/TimeStampValue[22]\, B
         => \MemorySynchronizer_0/TimeStampReg_Z[22]\, C => 
        ADLIB_GND0, D => ADLIB_GND0, FCI => 
        \MemorySynchronizer_0/temp_1_cry_21\, S => 
        \MemorySynchronizer_0/temp_1[22]\, Y => OPEN, FCO => 
        \MemorySynchronizer_0/temp_1_cry_22\, CC => 
        NET_CC_CONFIG265, P => NET_CC_CONFIG263, UB => 
        NET_CC_CONFIG264);
    
    \STAMP_0/un1_spi_rx_data_1[27]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame[59]\, B => 
        \STAMP_0/dummy_Z[27]\, C => \sb_sb_0_STAMP_PADDR[8]\, D
         => \sb_sb_0_STAMP_PADDR[9]\, Y => \STAMP_0/N_644\);
    
    \resetn_obuf/U0/U_IOPAD\ : sdf_IOPAD_TRI
      port map(PAD => resetn, D => \resetn_obuf/U0/DOUT\, E => 
        \resetn_obuf/U0/EOUT\);
    
    GND_power_inst1 : GND
      port map( Y => GND_power_net1);

    VCC_power_inst1 : VCC
      port map( Y => VCC_power_net1);


end DEF_ARCH; 
