-- ********************************************************************/
-- Actel Corporation Proprietary and Confidential
-- Copyright 2010 Actel Corporation.  All rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
-- ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
-- IN ADVANCE IN WRITING.
--
-- Description:         CoreAPB3 parameters
--
-- Revision Information:
-- Date			Description
-- ----			-----------------------------------------
-- 03Nov09		Production Release Version 3.0
--
-- SVN Revision Information:
-- SVN $Revision: 23124 $
-- SVN $Date: 2014-07-17 15:31:27 +0100 (Thu, 17 Jul 2014) $
--
-- Resolved SARs
-- SAR      Date     Who   Description
--
-- Notes:
--
-- *********************************************************************/

package coreparameters is
    constant APBSLOT0ENABLE : integer := 1;
    constant APBSLOT10ENABLE : integer := 1;
    constant APBSLOT11ENABLE : integer := 1;
    constant APBSLOT12ENABLE : integer := 1;
    constant APBSLOT13ENABLE : integer := 1;
    constant APBSLOT14ENABLE : integer := 1;
    constant APBSLOT15ENABLE : integer := 1;
    constant APBSLOT1ENABLE : integer := 1;
    constant APBSLOT2ENABLE : integer := 1;
    constant APBSLOT3ENABLE : integer := 1;
    constant APBSLOT4ENABLE : integer := 1;
    constant APBSLOT5ENABLE : integer := 1;
    constant APBSLOT6ENABLE : integer := 1;
    constant APBSLOT7ENABLE : integer := 1;
    constant APBSLOT8ENABLE : integer := 1;
    constant APBSLOT9ENABLE : integer := 1;
    constant APB_DWIDTH : integer := 32;
    constant IADDR_OPTION : integer := 0;
    constant MADDR_BITS : integer := 32;
    constant SC_0 : integer := 0;
    constant SC_1 : integer := 0;
    constant SC_10 : integer := 0;
    constant SC_11 : integer := 0;
    constant SC_12 : integer := 0;
    constant SC_13 : integer := 0;
    constant SC_14 : integer := 0;
    constant SC_15 : integer := 0;
    constant SC_2 : integer := 0;
    constant SC_3 : integer := 0;
    constant SC_4 : integer := 0;
    constant SC_5 : integer := 0;
    constant SC_6 : integer := 0;
    constant SC_7 : integer := 0;
    constant SC_8 : integer := 0;
    constant SC_9 : integer := 0;
    constant UPR_NIBBLE_POSN : integer := 7;
	constant FAMILY          : integer := 19;
end coreparameters;
