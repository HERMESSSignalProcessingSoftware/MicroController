-- Version: v12.6 12.900.20.24

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity spi_master_2_32 is

    port( SPITransmitReg    : in    std_logic_vector(31 downto 0);
          SPIaddr_0         : in    std_logic;
          SPIRecReg         : out   std_logic_vector(31 downto 0);
          enable            : in    std_logic;
          InternalBusy      : out   std_logic;
          mosi_cl_1z        : out   std_logic;
          mosi_1_1z         : out   std_logic;
          resetn            : in    std_logic;
          SCLK_c            : out   std_logic;
          MISO_c            : in    std_logic;
          nCS2_c            : out   std_logic;
          resetn_arst       : in    std_logic;
          nCS1_c            : out   std_logic;
          sb_sb_0_FIC_0_CLK : in    std_logic
        );

end spi_master_2_32;

architecture DEF_ARCH of spi_master_2_32 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \mosi_cl_1z\, \SCLK_c\, \nCS2_c\, \nCS1_c\
         : std_logic;
    signal rx_buffer_Z : std_logic_vector(31 downto 0);
    signal ss_n_buffer_5 : std_logic_vector(1 downto 0);
    signal tx_buffer_Z : std_logic_vector(31 downto 0);
    signal tx_buffer_RNO_Z : std_logic_vector(30 downto 0);
    signal slave_Z : std_logic_vector(0 to 0);
    signal state_Z : std_logic_vector(0 to 0);
    signal count_Z : std_logic_vector(31 downto 0);
    signal count_lm : std_logic_vector(31 downto 0);
    signal clk_toggles_Z : std_logic_vector(6 downto 0);
    signal clk_toggles_s : std_logic_vector(6 downto 0);
    signal clk_toggles_cry : std_logic_vector(5 downto 0);
    signal clk_toggles_RNIIG4O1_Y : std_logic_vector(0 to 0);
    signal clk_toggles_RNIFEQO2_Y : std_logic_vector(1 to 1);
    signal clk_toggles_RNIDDGP3_Y : std_logic_vector(2 to 2);
    signal clk_toggles_RNICD6Q4_Y : std_logic_vector(3 to 3);
    signal clk_toggles_RNICESQ5_Y : std_logic_vector(4 to 4);
    signal clk_toggles_RNO_FCO : std_logic_vector(6 to 6);
    signal clk_toggles_RNO_Y : std_logic_vector(6 to 6);
    signal clk_toggles_RNIDGIR6_Y : std_logic_vector(5 to 5);
    signal count_cry_Z : std_logic_vector(30 downto 1);
    signal count_s : std_logic_vector(30 downto 1);
    signal count_cry_Y_0 : std_logic_vector(30 downto 1);
    signal count_s_FCO_0 : std_logic_vector(31 to 31);
    signal count_s_Z : std_logic_vector(31 to 31);
    signal count_s_Y_0 : std_logic_vector(31 to 31);
    signal \VCC\, rx_buffer_0_sqmuxa_1, \GND\, 
        un1_reset_n_inv_2_i, N_4390, N_4402, N_4417, N_15_i, N_20, 
        assert_data_Z, N_18_i, mosi_1_3, count_0_sqmuxa, busy_15, 
        N_28_i, N_4_i, N_46, clk_toggles_cry_cy, 
        un10_count_0_a2_RNIMJEN_S, un10_count_0_a2_RNIMJEN_Y, 
        un10_count_i, count_s_834_FCO, count_s_834_S, 
        count_s_834_Y, un7_count_NE_i, un7_count_NE_13_Z, 
        un10_count_0_o2_0_Z, N_32, mosi_1_3_0_0_a2_0_Z, 
        un7_count_NE_23_Z, un7_count_NE_21_Z, un7_count_NE_20_Z, 
        un7_count_NE_19_Z, un7_count_NE_18_Z, un7_count_NE_17_Z, 
        un7_count_NE_16_Z, ss_n_buffer_1_sqmuxa_0_a2_Z, N_47, 
        un7_count_NE_27_Z, N_42, un7_count_NE_28_Z, N_13_i, N_45, 
        rx_buffer_0_sqmuxa_1_tz, N_1488, N_68, N_67 : std_logic;

begin 

    mosi_cl_1z <= \mosi_cl_1z\;
    SCLK_c <= \SCLK_c\;
    nCS2_c <= \nCS2_c\;
    nCS1_c <= \nCS1_c\;

    \tx_buffer[28]\ : SLE
      port map(D => tx_buffer_RNO_Z(28), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(28));
    
    \rx_buffer[16]\ : SLE
      port map(D => rx_buffer_Z(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(16));
    
    \count_lm_0[13]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(13), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(13));
    
    \count[27]\ : SLE
      port map(D => count_lm(27), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(27));
    
    \rx_buffer[11]\ : SLE
      port map(D => rx_buffer_Z(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(11));
    
    \state[0]\ : SLE
      port map(D => busy_15, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => state_Z(0));
    
    \count[25]\ : SLE
      port map(D => count_lm(25), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(25));
    
    \tx_buffer_RNO[14]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(14), B => state_Z(0), C => 
        tx_buffer_Z(13), Y => tx_buffer_RNO_Z(14));
    
    \count[17]\ : SLE
      port map(D => count_lm(17), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(17));
    
    un10_count_0_o2 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => clk_toggles_Z(1), B => un10_count_0_o2_0_Z, C
         => clk_toggles_Z(5), D => clk_toggles_Z(2), Y => N_42);
    
    \tx_buffer[16]\ : SLE
      port map(D => tx_buffer_RNO_Z(16), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(16));
    
    \tx_buffer[11]\ : SLE
      port map(D => tx_buffer_RNO_Z(11), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(11));
    
    \count[15]\ : SLE
      port map(D => count_lm(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(15));
    
    \tx_buffer_RNO[23]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(23), B => state_Z(0), C => 
        tx_buffer_Z(22), Y => tx_buffer_RNO_Z(23));
    
    rx_buffer_0_sqmuxa_1_0_tz : CFG4
      generic map(INIT => x"1050")

      port map(A => N_32, B => clk_toggles_Z(6), C => resetn, D
         => N_45, Y => rx_buffer_0_sqmuxa_1_tz);
    
    \rx_buffer[17]\ : SLE
      port map(D => rx_buffer_Z(16), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(17));
    
    \count_cry[14]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(14), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(13), S => count_s(14), Y => 
        count_cry_Y_0(14), FCO => count_cry_Z(14));
    
    \rx_data[2]\ : SLE
      port map(D => rx_buffer_Z(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(2));
    
    sclk_buffer_0_sqmuxa_i_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => N_42, B => clk_toggles_Z(0), Y => N_45);
    
    \tx_buffer[17]\ : SLE
      port map(D => N_4417, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(17));
    
    \count[9]\ : SLE
      port map(D => count_lm(9), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(9));
    
    \tx_buffer[29]\ : SLE
      port map(D => tx_buffer_RNO_Z(29), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(29));
    
    \rx_data[30]\ : SLE
      port map(D => rx_buffer_Z(30), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(30));
    
    sclk_buffer_6_iv_i_0_RNO : CFG4
      generic map(INIT => x"1050")

      port map(A => N_32, B => clk_toggles_Z(6), C => 
        un7_count_NE_i, D => N_45, Y => N_13_i);
    
    \count_lm_0[17]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(17), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(17));
    
    \rx_data[21]\ : SLE
      port map(D => rx_buffer_Z(21), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(21));
    
    \tx_buffer_RNO[30]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(30), B => state_Z(0), C => 
        tx_buffer_Z(29), Y => tx_buffer_RNO_Z(30));
    
    \rx_buffer[20]\ : SLE
      port map(D => rx_buffer_Z(19), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(20));
    
    \count_cry[28]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(28), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(27), S => count_s(28), Y => 
        count_cry_Y_0(28), FCO => count_cry_Z(28));
    
    \count[8]\ : SLE
      port map(D => count_lm(8), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(8));
    
    \count_cry[26]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(26), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(25), S => count_s(26), Y => 
        count_cry_Y_0(26), FCO => count_cry_Z(26));
    
    \rx_data[16]\ : SLE
      port map(D => rx_buffer_Z(16), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(16));
    
    \rx_data[15]\ : SLE
      port map(D => rx_buffer_Z(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(15));
    
    \count_cry[20]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(20), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(19), S => count_s(20), Y => 
        count_cry_Y_0(20), FCO => count_cry_Z(20));
    
    \count_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(8), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(7), S => count_s(8), Y => 
        count_cry_Y_0(8), FCO => count_cry_Z(8));
    
    \count_lm_0[6]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(6), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(6));
    
    \rx_data[3]\ : SLE
      port map(D => rx_buffer_Z(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(3));
    
    \tx_buffer_RNO[25]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(25), B => state_Z(0), C => 
        tx_buffer_Z(24), Y => tx_buffer_RNO_Z(25));
    
    \rx_data[7]\ : SLE
      port map(D => rx_buffer_Z(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(7));
    
    \tx_buffer[5]\ : SLE
      port map(D => tx_buffer_RNO_Z(5), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(5));
    
    \tx_buffer_RNO[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(1), B => state_Z(0), C => 
        tx_buffer_Z(0), Y => tx_buffer_RNO_Z(1));
    
    \rx_buffer[24]\ : SLE
      port map(D => rx_buffer_Z(23), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(24));
    
    \tx_buffer_RNO[13]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(13), B => state_Z(0), C => 
        tx_buffer_Z(12), Y => tx_buffer_RNO_Z(13));
    
    \rx_buffer[10]\ : SLE
      port map(D => rx_buffer_Z(9), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(10));
    
    \count[20]\ : SLE
      port map(D => count_lm(20), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(20));
    
    \rx_data[4]\ : SLE
      port map(D => rx_buffer_Z(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(4));
    
    \tx_buffer[10]\ : SLE
      port map(D => tx_buffer_RNO_Z(10), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(10));
    
    \count_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(2), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(1), S => count_s(2), Y => 
        count_cry_Y_0(2), FCO => count_cry_Z(2));
    
    \count[10]\ : SLE
      port map(D => count_lm(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(10));
    
    \tx_buffer[7]\ : SLE
      port map(D => tx_buffer_RNO_Z(7), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(7));
    
    \tx_buffer[3]\ : SLE
      port map(D => tx_buffer_RNO_Z(3), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(3));
    
    \rx_buffer[23]\ : SLE
      port map(D => rx_buffer_Z(22), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(23));
    
    \count_lm_0[5]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(5), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(5));
    
    \count_lm_0[28]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(28), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(28));
    
    \count_cry[15]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(15), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(14), S => count_s(15), Y => 
        count_cry_Y_0(15), FCO => count_cry_Z(15));
    
    \count[5]\ : SLE
      port map(D => count_lm(5), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(5));
    
    un10_count_0_a2_RNIMJEN : ARI1
      generic map(INIT => x"42200")

      port map(A => \VCC\, B => state_Z(0), C => un10_count_i, D
         => \GND\, FCI => \VCC\, S => un10_count_0_a2_RNIMJEN_S, 
        Y => un10_count_0_a2_RNIMJEN_Y, FCO => clk_toggles_cry_cy);
    
    \rx_buffer[14]\ : SLE
      port map(D => rx_buffer_Z(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(14));
    
    ss_n_buffer_1_sqmuxa_0_a2 : CFG3
      generic map(INIT => x"4C")

      port map(A => un7_count_NE_i, B => state_Z(0), C => 
        un10_count_i, Y => ss_n_buffer_1_sqmuxa_0_a2_Z);
    
    \tx_buffer_RNO[9]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(9), B => state_Z(0), C => 
        tx_buffer_Z(8), Y => tx_buffer_RNO_Z(9));
    
    \count_s[31]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(31), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(30), S => count_s_Z(31), Y => 
        count_s_Y_0(31), FCO => count_s_FCO_0(31));
    
    \tx_buffer_RNO[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(6), B => state_Z(0), C => 
        tx_buffer_Z(5), Y => tx_buffer_RNO_Z(6));
    
    \tx_buffer[14]\ : SLE
      port map(D => tx_buffer_RNO_Z(14), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(14));
    
    \rx_data[5]\ : SLE
      port map(D => rx_buffer_Z(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(5));
    
    \rx_buffer[7]\ : SLE
      port map(D => rx_buffer_Z(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(7));
    
    count_s_834 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(0), C => \GND\, D => 
        \GND\, FCI => \VCC\, S => count_s_834_S, Y => 
        count_s_834_Y, FCO => count_s_834_FCO);
    
    \rx_buffer[13]\ : SLE
      port map(D => rx_buffer_Z(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(13));
    
    un7_count_NE_16 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(4), B => count_Z(3), C => count_Z(1), 
        D => count_Z(0), Y => un7_count_NE_16_Z);
    
    \state_RNIS9IF2[0]\ : CFG4
      generic map(INIT => x"E200")

      port map(A => enable, B => state_Z(0), C => un7_count_NE_i, 
        D => resetn, Y => N_46);
    
    \clk_toggles_RNICESQ5[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => un10_count_0_a2_RNIMJEN_Y, C => 
        clk_toggles_Z(4), D => \GND\, FCI => clk_toggles_cry(3), 
        S => clk_toggles_s(4), Y => clk_toggles_RNICESQ5_Y(4), 
        FCO => clk_toggles_cry(4));
    
    \tx_buffer_RNO[15]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(15), B => state_Z(0), C => 
        tx_buffer_Z(14), Y => tx_buffer_RNO_Z(15));
    
    \count_cry[30]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(30), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(29), S => count_s(30), Y => 
        count_cry_Y_0(30), FCO => count_cry_Z(30));
    
    \count_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(12), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(11), S => count_s(12), Y => 
        count_cry_Y_0(12), FCO => count_cry_Z(12));
    
    \tx_buffer_RNO[27]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(27), B => state_Z(0), C => 
        tx_buffer_Z(26), Y => tx_buffer_RNO_Z(27));
    
    \tx_buffer[13]\ : SLE
      port map(D => tx_buffer_RNO_Z(13), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(13));
    
    \count_lm_0[24]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(24), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(24));
    
    \count_cry[19]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(19), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(18), S => count_s(19), Y => 
        count_cry_Y_0(19), FCO => count_cry_Z(19));
    
    \count[4]\ : SLE
      port map(D => count_lm(4), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(4));
    
    un10_count_0_a2_RNIQST32 : CFG3
      generic map(INIT => x"80")

      port map(A => un7_count_NE_i, B => state_Z(0), C => 
        un10_count_i, Y => N_15_i);
    
    sclk_buffer_0_sqmuxa_i_0_m2 : CFG3
      generic map(INIT => x"E2")

      port map(A => \nCS1_c\, B => slave_Z(0), C => \nCS2_c\, Y
         => N_32);
    
    \count[22]\ : SLE
      port map(D => count_lm(22), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(22));
    
    \rx_data[24]\ : SLE
      port map(D => rx_buffer_Z(24), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(24));
    
    mosi_1 : SLE
      port map(D => tx_buffer_Z(31), CLK => sb_sb_0_FIC_0_CLK, EN
         => mosi_1_3, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => mosi_1_1z);
    
    \count[12]\ : SLE
      port map(D => count_lm(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(12));
    
    \state_RNIO0331[0]\ : CFG3
      generic map(INIT => x"E0")

      port map(A => enable, B => state_Z(0), C => resetn, Y => 
        N_4_i);
    
    \count_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(6), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(5), S => count_s(6), Y => 
        count_cry_Y_0(6), FCO => count_cry_Z(6));
    
    \count[0]\ : SLE
      port map(D => count_lm(0), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(0));
    
    assert_data_RNO : CFG4
      generic map(INIT => x"52A2")

      port map(A => assert_data_Z, B => enable, C => state_Z(0), 
        D => un7_count_NE_i, Y => N_18_i);
    
    \rx_data[11]\ : SLE
      port map(D => rx_buffer_Z(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(11));
    
    \tx_buffer_RNO[31]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(31), B => state_Z(0), C => 
        tx_buffer_Z(30), Y => N_4402);
    
    \count_lm_0[21]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(21), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(21));
    
    \count_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(5), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(4), S => count_s(5), Y => 
        count_cry_Y_0(5), FCO => count_cry_Z(5));
    
    \tx_buffer[26]\ : SLE
      port map(D => tx_buffer_RNO_Z(26), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(26));
    
    \tx_buffer[21]\ : SLE
      port map(D => tx_buffer_RNO_Z(21), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(21));
    
    \tx_buffer_RNO[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(2), B => state_Z(0), C => 
        tx_buffer_Z(1), Y => tx_buffer_RNO_Z(2));
    
    rx_buffer_0_sqmuxa_1_0 : CFG4
      generic map(INIT => x"2000")

      port map(A => state_Z(0), B => assert_data_Z, C => 
        rx_buffer_0_sqmuxa_1_tz, D => un7_count_NE_i, Y => 
        rx_buffer_0_sqmuxa_1);
    
    \tx_buffer_RNO[17]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(17), B => state_Z(0), C => 
        tx_buffer_Z(16), Y => N_4417);
    
    \rx_buffer[8]\ : SLE
      port map(D => rx_buffer_Z(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(8));
    
    \tx_buffer[27]\ : SLE
      port map(D => tx_buffer_RNO_Z(27), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(27));
    
    \tx_buffer[9]\ : SLE
      port map(D => tx_buffer_RNO_Z(9), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(9));
    
    \count_lm_0[8]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(8), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(8));
    
    \tx_buffer_RNO[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(4), B => state_Z(0), C => 
        tx_buffer_Z(3), Y => tx_buffer_RNO_Z(4));
    
    \tx_buffer[2]\ : SLE
      port map(D => tx_buffer_RNO_Z(2), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(2));
    
    \count_lm_0[10]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(10), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(10));
    
    \rx_buffer[5]\ : SLE
      port map(D => rx_buffer_Z(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(5));
    
    count_0_sqmuxa_0_a2 : CFG3
      generic map(INIT => x"20")

      port map(A => enable, B => state_Z(0), C => resetn, Y => 
        count_0_sqmuxa);
    
    \count_lm_0[29]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(29), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(29));
    
    \rx_buffer[4]\ : SLE
      port map(D => rx_buffer_Z(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(4));
    
    \count_cry[21]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(21), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(20), S => count_s(21), Y => 
        count_cry_Y_0(21), FCO => count_cry_Z(21));
    
    \count[23]\ : SLE
      port map(D => count_lm(23), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(23));
    
    busy : SLE
      port map(D => busy_15, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \GND\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => InternalBusy);
    
    \count[13]\ : SLE
      port map(D => count_lm(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(13));
    
    \tx_buffer_RNO[28]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(28), B => state_Z(0), C => 
        tx_buffer_Z(27), Y => tx_buffer_RNO_Z(28));
    
    \count_cry[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(13), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(12), S => count_s(13), Y => 
        count_cry_Y_0(13), FCO => count_cry_Z(13));
    
    \count_cry[24]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(24), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(23), S => count_s(24), Y => 
        count_cry_Y_0(24), FCO => count_cry_Z(24));
    
    \count_cry[17]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(17), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(16), S => count_s(17), Y => 
        count_cry_Y_0(17), FCO => count_cry_Z(17));
    
    GND_Z : GND
      port map(Y => \GND\);
    
    un7_count_NE_17 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(8), B => count_Z(7), C => count_Z(6), 
        D => count_Z(5), Y => un7_count_NE_17_Z);
    
    un10_count_0_a2 : CFG3
      generic map(INIT => x"20")

      port map(A => clk_toggles_Z(6), B => N_42, C => 
        clk_toggles_Z(0), Y => un10_count_i);
    
    \rx_buffer[25]\ : SLE
      port map(D => rx_buffer_Z(24), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(25));
    
    un7_count_NE_18 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(12), B => count_Z(11), C => 
        count_Z(10), D => count_Z(9), Y => un7_count_NE_18_Z);
    
    \rx_buffer[22]\ : SLE
      port map(D => rx_buffer_Z(21), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(22));
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    \tx_buffer[20]\ : SLE
      port map(D => tx_buffer_RNO_Z(20), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(20));
    
    \count_lm_0[0]\ : CFG4
      generic map(INIT => x"2733")

      port map(A => un7_count_NE_i, B => count_0_sqmuxa, C => 
        count_Z(0), D => state_Z(0), Y => count_lm(0));
    
    \count_lm_0[25]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(25), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(25));
    
    un7_count_NE_13 : CFG2
      generic map(INIT => x"E")

      port map(A => count_Z(27), B => count_Z(28), Y => 
        un7_count_NE_13_Z);
    
    \rx_data[1]\ : SLE
      port map(D => rx_buffer_Z(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(1));
    
    \rx_buffer[1]\ : SLE
      port map(D => rx_buffer_Z(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(1));
    
    \rx_data[14]\ : SLE
      port map(D => rx_buffer_Z(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(14));
    
    \count[1]\ : SLE
      port map(D => count_lm(1), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(1));
    
    \clk_toggles_RNO[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => un10_count_0_a2_RNIMJEN_Y, C => 
        clk_toggles_Z(6), D => \GND\, FCI => clk_toggles_cry(5), 
        S => clk_toggles_s(6), Y => clk_toggles_RNO_Y(6), FCO => 
        clk_toggles_RNO_FCO(6));
    
    \count[3]\ : SLE
      port map(D => count_lm(3), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(3));
    
    \tx_buffer[24]\ : SLE
      port map(D => tx_buffer_RNO_Z(24), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(24));
    
    \rx_data[20]\ : SLE
      port map(D => rx_buffer_Z(20), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(20));
    
    \rx_buffer[15]\ : SLE
      port map(D => rx_buffer_Z(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(15));
    
    \clk_toggles[2]\ : SLE
      port map(D => clk_toggles_s(2), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_46, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => clk_toggles_Z(2));
    
    \rx_data[22]\ : SLE
      port map(D => rx_buffer_Z(22), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(22));
    
    \rx_buffer[12]\ : SLE
      port map(D => rx_buffer_Z(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(12));
    
    \count_lm_0[4]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(4), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(4));
    
    \count_lm_0[22]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(22), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(22));
    
    \count[29]\ : SLE
      port map(D => count_lm(29), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(29));
    
    \count_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(7), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(6), S => count_s(7), Y => 
        count_cry_Y_0(7), FCO => count_cry_Z(7));
    
    \tx_buffer[15]\ : SLE
      port map(D => tx_buffer_RNO_Z(15), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(15));
    
    \count[19]\ : SLE
      port map(D => count_lm(19), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(19));
    
    \tx_buffer[12]\ : SLE
      port map(D => tx_buffer_RNO_Z(12), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(12));
    
    \rx_data[28]\ : SLE
      port map(D => rx_buffer_Z(28), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(28));
    
    \tx_buffer_RNO[18]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(18), B => state_Z(0), C => 
        tx_buffer_Z(17), Y => tx_buffer_RNO_Z(18));
    
    \ss_n_buffer_5_0[0]\ : CFG3
      generic map(INIT => x"B3")

      port map(A => \nCS1_c\, B => ss_n_buffer_1_sqmuxa_0_a2_Z, C
         => slave_Z(0), Y => ss_n_buffer_5(0));
    
    \count_lm_0[18]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(18), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(18));
    
    un7_count_NE_27 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(25), B => count_Z(26), C => 
        un7_count_NE_23_Z, D => un7_count_NE_13_Z, Y => 
        un7_count_NE_27_Z);
    
    un7_count_NE_28 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un7_count_NE_19_Z, B => un7_count_NE_18_Z, C
         => un7_count_NE_17_Z, D => un7_count_NE_16_Z, Y => 
        un7_count_NE_28_Z);
    
    \tx_buffer[23]\ : SLE
      port map(D => tx_buffer_RNO_Z(23), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(23));
    
    sclk_buffer_6_iv_i_0 : CFG4
      generic map(INIT => x"33D8")

      port map(A => state_Z(0), B => N_13_i, C => enable, D => 
        \SCLK_c\, Y => N_20);
    
    \clk_toggles[0]\ : SLE
      port map(D => clk_toggles_s(0), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_46, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => clk_toggles_Z(0));
    
    \tx_buffer[4]\ : SLE
      port map(D => tx_buffer_RNO_Z(4), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(4));
    
    \count_lm_0[30]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(30), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(30));
    
    un7_count_NE_23 : CFG4
      generic map(INIT => x"FEFF")

      port map(A => count_Z(31), B => count_Z(30), C => 
        count_Z(29), D => count_Z(2), Y => un7_count_NE_23_Z);
    
    \tx_buffer[31]\ : SLE
      port map(D => N_4402, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(31));
    
    \count_cry[25]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(25), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(24), S => count_s(25), Y => 
        count_cry_Y_0(25), FCO => count_cry_Z(25));
    
    \clk_toggles[1]\ : SLE
      port map(D => clk_toggles_s(1), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_46, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => clk_toggles_Z(1));
    
    un7_count_NE_20_RNI49FC1 : CFG4
      generic map(INIT => x"0001")

      port map(A => un7_count_NE_20_Z, B => un7_count_NE_21_Z, C
         => un7_count_NE_28_Z, D => un7_count_NE_27_Z, Y => 
        un7_count_NE_i);
    
    sclk_buffer : SLE
      port map(D => N_20, CLK => sb_sb_0_FIC_0_CLK, EN => resetn, 
        ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => \GND\, 
        LAT => \GND\, Q => \SCLK_c\);
    
    \count_lm_0[26]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(26), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(26));
    
    \count_lm_0[9]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(9), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(9));
    
    \rx_buffer[3]\ : SLE
      port map(D => rx_buffer_Z(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(3));
    
    \tx_buffer[8]\ : SLE
      port map(D => tx_buffer_RNO_Z(8), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(8));
    
    \rx_data[29]\ : SLE
      port map(D => rx_buffer_Z(29), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(29));
    
    \count_lm_0[14]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(14), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(14));
    
    un7_count_NE_19 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(16), B => count_Z(15), C => 
        count_Z(14), D => count_Z(13), Y => un7_count_NE_19_Z);
    
    \tx_buffer_RNO[22]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(22), B => state_Z(0), C => 
        tx_buffer_Z(21), Y => tx_buffer_RNO_Z(22));
    
    \tx_buffer[6]\ : SLE
      port map(D => tx_buffer_RNO_Z(6), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(6));
    
    \count_cry[22]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(22), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(21), S => count_s(22), Y => 
        count_cry_Y_0(22), FCO => count_cry_Z(22));
    
    \count_cry[29]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(29), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(28), S => count_s(29), Y => 
        count_cry_Y_0(29), FCO => count_cry_Z(29));
    
    \tx_buffer_RNO[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => state_Z(0), B => SPITransmitReg(0), Y => 
        tx_buffer_RNO_Z(0));
    
    un7_count_NE_20 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(20), B => count_Z(19), C => 
        count_Z(18), D => count_Z(17), Y => un7_count_NE_20_Z);
    
    \rx_buffer[28]\ : SLE
      port map(D => rx_buffer_Z(27), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(28));
    
    \rx_data[31]\ : SLE
      port map(D => rx_buffer_Z(31), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(31));
    
    \tx_buffer_RNO[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(5), B => state_Z(0), C => 
        tx_buffer_Z(4), Y => tx_buffer_RNO_Z(5));
    
    \count_lm_0[23]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(23), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(23));
    
    \count_lm_0[1]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(1), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(1));
    
    \rx_buffer[6]\ : SLE
      port map(D => rx_buffer_Z(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(6));
    
    \clk_toggles_RNIIG4O1[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => un10_count_0_a2_RNIMJEN_Y, C => 
        clk_toggles_Z(0), D => \GND\, FCI => clk_toggles_cry_cy, 
        S => clk_toggles_s(0), Y => clk_toggles_RNIIG4O1_Y(0), 
        FCO => clk_toggles_cry(0));
    
    \tx_buffer_RNO[20]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(20), B => state_Z(0), C => 
        tx_buffer_Z(19), Y => tx_buffer_RNO_Z(20));
    
    \clk_toggles_RNICD6Q4[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => un10_count_0_a2_RNIMJEN_Y, C => 
        clk_toggles_Z(3), D => \GND\, FCI => clk_toggles_cry(2), 
        S => clk_toggles_s(3), Y => clk_toggles_RNICD6Q4_Y(3), 
        FCO => clk_toggles_cry(3));
    
    \slave[0]\ : SLE
      port map(D => SPIaddr_0, CLK => sb_sb_0_FIC_0_CLK, EN => 
        count_0_sqmuxa, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => slave_Z(0));
    
    \rx_buffer[29]\ : SLE
      port map(D => rx_buffer_Z(28), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(29));
    
    un10_count_0_o2_0 : CFG2
      generic map(INIT => x"E")

      port map(A => clk_toggles_Z(3), B => clk_toggles_Z(4), Y
         => un10_count_0_o2_0_Z);
    
    \clk_toggles[4]\ : SLE
      port map(D => clk_toggles_s(4), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_46, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => clk_toggles_Z(4));
    
    \count_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(4), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(3), S => count_s(4), Y => 
        count_cry_Y_0(4), FCO => count_cry_Z(4));
    
    \count_lm_0[11]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(11), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(11));
    
    \rx_data[23]\ : SLE
      port map(D => rx_buffer_Z(23), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(23));
    
    \clk_toggles_RNIDGIR6[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => un10_count_0_a2_RNIMJEN_Y, C => 
        clk_toggles_Z(5), D => \GND\, FCI => clk_toggles_cry(4), 
        S => clk_toggles_s(5), Y => clk_toggles_RNIDGIR6_Y(5), 
        FCO => clk_toggles_cry(5));
    
    \tx_buffer[30]\ : SLE
      port map(D => tx_buffer_RNO_Z(30), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(30));
    
    \rx_buffer[31]\ : SLE
      port map(D => rx_buffer_Z(30), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(31));
    
    \rx_buffer[18]\ : SLE
      port map(D => rx_buffer_Z(17), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(18));
    
    \count_cry[18]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(18), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(17), S => count_s(18), Y => 
        count_cry_Y_0(18), FCO => count_cry_Z(18));
    
    \count_lm_0[27]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(27), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(27));
    
    \count_cry[16]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(16), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(15), S => count_s(16), Y => 
        count_cry_Y_0(16), FCO => count_cry_Z(16));
    
    \tx_buffer[1]\ : SLE
      port map(D => tx_buffer_RNO_Z(1), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(1));
    
    \tx_buffer[18]\ : SLE
      port map(D => tx_buffer_RNO_Z(18), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(18));
    
    \rx_buffer[2]\ : SLE
      port map(D => rx_buffer_Z(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(2));
    
    \count_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(10), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(9), S => count_s(10), Y => 
        count_cry_Y_0(10), FCO => count_cry_Z(10));
    
    \tx_buffer_RNO[12]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(12), B => state_Z(0), C => 
        tx_buffer_Z(11), Y => tx_buffer_RNO_Z(12));
    
    \rx_data[10]\ : SLE
      port map(D => rx_buffer_Z(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(10));
    
    \rx_data[12]\ : SLE
      port map(D => rx_buffer_Z(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(12));
    
    \rx_buffer[19]\ : SLE
      port map(D => rx_buffer_Z(18), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(19));
    
    \count[31]\ : SLE
      port map(D => count_lm(31), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(31));
    
    \rx_data[27]\ : SLE
      port map(D => rx_buffer_Z(27), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(27));
    
    \count[28]\ : SLE
      port map(D => count_lm(28), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(28));
    
    mosi_1_3_0_0_a2_0 : CFG3
      generic map(INIT => x"20")

      port map(A => assert_data_Z, B => clk_toggles_Z(6), C => 
        resetn, Y => mosi_1_3_0_0_a2_0_Z);
    
    \tx_buffer[19]\ : SLE
      port map(D => N_4390, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(19));
    
    \rx_data[18]\ : SLE
      port map(D => rx_buffer_Z(18), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(18));
    
    \count_lm_0[19]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(19), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(19));
    
    \count[18]\ : SLE
      port map(D => count_lm(18), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(18));
    
    \count[7]\ : SLE
      port map(D => count_lm(7), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(7));
    
    \count_lm_0[3]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(3), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(3));
    
    \tx_buffer_RNO[10]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(10), B => state_Z(0), C => 
        tx_buffer_Z(9), Y => tx_buffer_RNO_Z(10));
    
    \tx_buffer_RNO[26]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(26), B => state_Z(0), C => 
        tx_buffer_Z(25), Y => tx_buffer_RNO_Z(26));
    
    \rx_buffer[0]\ : SLE
      port map(D => MISO_c, CLK => sb_sb_0_FIC_0_CLK, EN => 
        rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(0));
    
    \rx_buffer[9]\ : SLE
      port map(D => rx_buffer_Z(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(9));
    
    busy_15_0_0 : CFG4
      generic map(INIT => x"77F0")

      port map(A => un10_count_i, B => un7_count_NE_i, C => 
        enable, D => state_Z(0), Y => busy_15);
    
    \rx_data[8]\ : SLE
      port map(D => rx_buffer_Z(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(8));
    
    \count[6]\ : SLE
      port map(D => count_lm(6), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(6));
    
    \tx_buffer_RNO[29]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(29), B => state_Z(0), C => 
        tx_buffer_Z(28), Y => tx_buffer_RNO_Z(29));
    
    \rx_data[6]\ : SLE
      port map(D => rx_buffer_Z(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(6));
    
    \count_cry[23]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(23), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(22), S => count_s(23), Y => 
        count_cry_Y_0(23), FCO => count_cry_Z(23));
    
    \rx_data[19]\ : SLE
      port map(D => rx_buffer_Z(19), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(19));
    
    \rx_buffer[30]\ : SLE
      port map(D => rx_buffer_Z(29), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(30));
    
    \tx_buffer[25]\ : SLE
      port map(D => tx_buffer_RNO_Z(25), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(25));
    
    \tx_buffer[22]\ : SLE
      port map(D => tx_buffer_RNO_Z(22), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(22));
    
    \ss_n_buffer[0]\ : SLE
      port map(D => ss_n_buffer_5(0), CLK => sb_sb_0_FIC_0_CLK, 
        EN => \VCC\, ALn => resetn_arst, ADn => \GND\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => \nCS1_c\);
    
    mosi_1_3_0_0_a2 : CFG4
      generic map(INIT => x"4000")

      port map(A => un10_count_i, B => state_Z(0), C => 
        mosi_1_3_0_0_a2_0_Z, D => un7_count_NE_i, Y => mosi_1_3);
    
    \count_cry[27]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(27), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(26), S => count_s(27), Y => 
        count_cry_Y_0(27), FCO => count_cry_Z(27));
    
    \count_lm_0[15]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(15), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(15));
    
    \rx_data[0]\ : SLE
      port map(D => rx_buffer_Z(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(0));
    
    assert_data_RNISDFD3 : CFG4
      generic map(INIT => x"44C4")

      port map(A => state_Z(0), B => N_46, C => assert_data_Z, D
         => clk_toggles_Z(6), Y => un1_reset_n_inv_2_i);
    
    \count[26]\ : SLE
      port map(D => count_lm(26), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(26));
    
    \tx_buffer[0]\ : SLE
      port map(D => tx_buffer_RNO_Z(0), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tx_buffer_Z(0));
    
    \count[16]\ : SLE
      port map(D => count_lm(16), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(16));
    
    \count_lm_0[31]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s_Z(31), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(31));
    
    \tx_buffer_RNO[8]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(8), B => state_Z(0), C => 
        tx_buffer_Z(7), Y => tx_buffer_RNO_Z(8));
    
    \count_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(3), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(2), S => count_s(3), Y => 
        count_cry_Y_0(3), FCO => count_cry_Z(3));
    
    \count[2]\ : SLE
      port map(D => count_lm(2), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(2));
    
    \clk_toggles[5]\ : SLE
      port map(D => clk_toggles_s(5), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_46, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => clk_toggles_Z(5));
    
    \tx_buffer_RNO[16]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(16), B => state_Z(0), C => 
        tx_buffer_Z(15), Y => tx_buffer_RNO_Z(16));
    
    \count_lm_0[12]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(12), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(12));
    
    \tx_buffer_RNO[21]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(21), B => state_Z(0), C => 
        tx_buffer_Z(20), Y => tx_buffer_RNO_Z(21));
    
    \clk_toggles_RNIDDGP3[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => un10_count_0_a2_RNIMJEN_Y, C => 
        clk_toggles_Z(2), D => \GND\, FCI => clk_toggles_cry(1), 
        S => clk_toggles_s(2), Y => clk_toggles_RNIDDGP3_Y(2), 
        FCO => clk_toggles_cry(2));
    
    \rx_data[26]\ : SLE
      port map(D => rx_buffer_Z(26), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(26));
    
    \rx_data[25]\ : SLE
      port map(D => rx_buffer_Z(25), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(25));
    
    \clk_toggles[3]\ : SLE
      port map(D => clk_toggles_s(3), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_46, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => clk_toggles_Z(3));
    
    un7_count_NE_21 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(24), B => count_Z(23), C => 
        count_Z(22), D => count_Z(21), Y => un7_count_NE_21_Z);
    
    \rx_data[13]\ : SLE
      port map(D => rx_buffer_Z(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(13));
    
    \tx_buffer_RNO[19]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(19), B => state_Z(0), C => 
        tx_buffer_Z(18), Y => N_4390);
    
    \tx_buffer_RNO[24]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(24), B => state_Z(0), C => 
        tx_buffer_Z(23), Y => tx_buffer_RNO_Z(24));
    
    \count[21]\ : SLE
      port map(D => count_lm(21), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(21));
    
    mosi_cl : SLE
      port map(D => N_28_i, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \mosi_cl_1z\);
    
    \count[11]\ : SLE
      port map(D => count_lm(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(11));
    
    \clk_toggles[6]\ : SLE
      port map(D => clk_toggles_s(6), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_46, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => clk_toggles_Z(6));
    
    \count_lm_0[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(7), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(7));
    
    \count_lm_0[2]\ : CFG4
      generic map(INIT => x"D8CC")

      port map(A => un7_count_NE_i, B => count_0_sqmuxa, C => 
        count_s(2), D => state_Z(0), Y => count_lm(2));
    
    \clk_toggles_RNIFEQO2[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => un10_count_0_a2_RNIMJEN_Y, C => 
        clk_toggles_Z(1), D => \GND\, FCI => clk_toggles_cry(0), 
        S => clk_toggles_s(1), Y => clk_toggles_RNIFEQO2_Y(1), 
        FCO => clk_toggles_cry(1));
    
    \count[24]\ : SLE
      port map(D => count_lm(24), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(24));
    
    \count[14]\ : SLE
      port map(D => count_lm(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(14));
    
    \rx_data[17]\ : SLE
      port map(D => rx_buffer_Z(17), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(17));
    
    \count_lm_0[16]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(16), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(16));
    
    \tx_buffer_RNO[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(7), B => state_Z(0), C => 
        tx_buffer_Z(6), Y => tx_buffer_RNO_Z(7));
    
    \rx_buffer[26]\ : SLE
      port map(D => rx_buffer_Z(25), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(26));
    
    \rx_buffer[21]\ : SLE
      port map(D => rx_buffer_Z(20), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(21));
    
    \rx_data[9]\ : SLE
      port map(D => rx_buffer_Z(9), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_15_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => SPIRecReg(9));
    
    \ss_n_buffer[1]\ : SLE
      port map(D => ss_n_buffer_5(1), CLK => sb_sb_0_FIC_0_CLK, 
        EN => \VCC\, ALn => resetn_arst, ADn => \GND\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => \nCS2_c\);
    
    \count[30]\ : SLE
      port map(D => count_lm(30), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_4_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(30));
    
    \ss_n_buffer_5_0[1]\ : CFG3
      generic map(INIT => x"3B")

      port map(A => \nCS2_c\, B => ss_n_buffer_1_sqmuxa_0_a2_Z, C
         => slave_Z(0), Y => ss_n_buffer_5(1));
    
    \tx_buffer_RNO[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(3), B => state_Z(0), C => 
        tx_buffer_Z(2), Y => tx_buffer_RNO_Z(3));
    
    \rx_buffer[27]\ : SLE
      port map(D => rx_buffer_Z(26), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(27));
    
    mosi_cl_RNO : CFG4
      generic map(INIT => x"D000")

      port map(A => N_47, B => \mosi_cl_1z\, C => resetn, D => 
        ss_n_buffer_1_sqmuxa_0_a2_Z, Y => N_28_i);
    
    assert_data : SLE
      port map(D => N_18_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        resetn, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => assert_data_Z);
    
    \tx_buffer_RNO[11]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => SPITransmitReg(11), B => state_Z(0), C => 
        tx_buffer_Z(10), Y => tx_buffer_RNO_Z(11));
    
    \count_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(11), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(10), S => count_s(11), Y => 
        count_cry_Y_0(11), FCO => count_cry_Z(11));
    
    \count_lm_0[20]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(20), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(20));
    
    \count_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(1), C => \GND\, D => 
        \GND\, FCI => count_s_834_FCO, S => count_s(1), Y => 
        count_cry_Y_0(1), FCO => count_cry_Z(1));
    
    mosi_cl_4_i_o2_0 : CFG3
      generic map(INIT => x"DF")

      port map(A => assert_data_Z, B => clk_toggles_Z(6), C => 
        un7_count_NE_i, Y => N_47);
    
    \count_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(9), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(8), S => count_s(9), Y => 
        count_cry_Y_0(9), FCO => count_cry_Z(9));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ram is

    port( InternalData2Memory : in    std_logic_vector(31 downto 0);
          InternalAddr2Memory : in    std_logic_vector(8 downto 0);
          InternalDataFromMem : out   std_logic_vector(31 downto 0);
          resetn              : in    std_logic;
          WriteEnable         : in    std_logic;
          sb_sb_0_FIC_0_CLK   : in    std_logic;
          resetn_arst         : in    std_logic
        );

end ram;

architecture DEF_ARCH of ram is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := ""; RAMINDEX:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \InternalDataFromMem\ : 
        std_logic_vector(31 downto 0);
    signal memory_memory_0_0_OLDA_Z : 
        std_logic_vector(31 downto 0);
    signal memory_memory_0_0_NEWA : 
        std_logic_vector(31 downto 0);
    signal memory_memory_0_0_A_DOUT : 
        std_logic_vector(17 downto 14);
    signal memoryro_507, \VCC\, memorywre_507, \GND\, 
        memoryro_508, memorywre_508, memoryro_509, memorywre_509, 
        memoryro_510, memorywre_510, memoryro_511, memorywre_511, 
        memoryro_502, memorywre_502, memoryro_503, memorywre_503, 
        memoryro_504, memorywre_504, memoryro_505, memorywre_505, 
        memoryro_506, memorywre_506, memoryro_497, memorywre_497, 
        memoryro_498, memorywre_498, memoryro_499, memorywre_499, 
        memoryro_500, memorywre_500, memoryro_501, memorywre_501, 
        memoryro_492, memorywre_492, memoryro_493, memorywre_493, 
        memoryro_494, memorywre_494, memoryro_495, memorywre_495, 
        memoryro_496, memorywre_496, memoryro_487, memorywre_487, 
        memoryro_488, memorywre_488, memoryro_489, memorywre_489, 
        memoryro_490, memorywre_490, memoryro_491, memorywre_491, 
        memoryro_482, memorywre_482, memoryro_483, memorywre_483, 
        memoryro_484, memorywre_484, memoryro_485, memorywre_485, 
        memoryro_486, memorywre_486, memoryro_477, memorywre_477, 
        memoryro_478, memorywre_478, memoryro_479, memorywre_479, 
        memoryro_480, memorywre_480, memoryro_481, memorywre_481, 
        memoryro_472, memorywre_472, memoryro_473, memorywre_473, 
        memoryro_474, memorywre_474, memoryro_475, memorywre_475, 
        memoryro_476, memorywre_476, memoryro_467, memorywre_467, 
        memoryro_468, memorywre_468, memoryro_469, memorywre_469, 
        memoryro_470, memorywre_470, memoryro_471, memorywre_471, 
        memoryro_462, memorywre_462, memoryro_463, memorywre_463, 
        memoryro_464, memorywre_464, memoryro_465, memorywre_465, 
        memoryro_466, memorywre_466, memoryro_457, memorywre_457, 
        memoryro_458, memorywre_458, memoryro_459, memorywre_459, 
        memoryro_460, memorywre_460, memoryro_461, memorywre_461, 
        memoryro_452, memorywre_452, memoryro_453, memorywre_453, 
        memoryro_454, memorywre_454, memoryro_455, memorywre_455, 
        memoryro_456, memorywre_456, memoryro_447, memorywre_447, 
        memoryro_448, memorywre_448, memoryro_449, memorywre_449, 
        memoryro_450, memorywre_450, memoryro_451, memorywre_451, 
        memoryro_442, memorywre_442, memoryro_443, memorywre_443, 
        memoryro_444, memorywre_444, memoryro_445, memorywre_445, 
        memoryro_446, memorywre_446, memoryro_437, memorywre_437, 
        memoryro_438, memorywre_438, memoryro_439, memorywre_439, 
        memoryro_440, memorywre_440, memoryro_441, memorywre_441, 
        memoryro_432, memorywre_432, memoryro_433, memorywre_433, 
        memoryro_434, memorywre_434, memoryro_435, memorywre_435, 
        memoryro_436, memorywre_436, memoryro_427, memorywre_427, 
        memoryro_428, memorywre_428, memoryro_429, memorywre_429, 
        memoryro_430, memorywre_430, memoryro_431, memorywre_431, 
        memoryro_422, memorywre_422, memoryro_423, memorywre_423, 
        memoryro_424, memorywre_424, memoryro_425, memorywre_425, 
        memoryro_426, memorywre_426, memoryro_417, memorywre_417, 
        memoryro_418, memorywre_418, memoryro_419, memorywre_419, 
        memoryro_420, memorywre_420, memoryro_421, memorywre_421, 
        memoryro_412, memorywre_412, memoryro_413, memorywre_413, 
        memoryro_414, memorywre_414, memoryro_415, memorywre_415, 
        memoryro_416, memorywre_416, memoryro_407, memorywre_407, 
        memoryro_408, memorywre_408, memoryro_409, memorywre_409, 
        memoryro_410, memorywre_410, memoryro_411, memorywre_411, 
        memoryro_402, memorywre_402, memoryro_403, memorywre_403, 
        memoryro_404, memorywre_404, memoryro_405, memorywre_405, 
        memoryro_406, memorywre_406, memoryro_397, memorywre_397, 
        memoryro_398, memorywre_398, memoryro_399, memorywre_399, 
        memoryro_400, memorywre_400, memoryro_401, memorywre_401, 
        memoryro_392, memorywre_392, memoryro_393, memorywre_393, 
        memoryro_394, memorywre_394, memoryro_395, memorywre_395, 
        memoryro_396, memorywre_396, memoryro_387, memorywre_387, 
        memoryro_388, memorywre_388, memoryro_389, memorywre_389, 
        memoryro_390, memorywre_390, memoryro_391, memorywre_391, 
        memoryro_382, memorywre_382, memoryro_383, memorywre_383, 
        memoryro_384, memorywre_384, memoryro_385, memorywre_385, 
        memoryro_386, memorywre_386, memoryro_377, memorywre_377, 
        memoryro_378, memorywre_378, memoryro_379, memorywre_379, 
        memoryro_380, memorywre_380, memoryro_381, memorywre_381, 
        memoryro_372, memorywre_372, memoryro_373, memorywre_373, 
        memoryro_374, memorywre_374, memoryro_375, memorywre_375, 
        memoryro_376, memorywre_376, memoryro_367, memorywre_367, 
        memoryro_368, memorywre_368, memoryro_369, memorywre_369, 
        memoryro_370, memorywre_370, memoryro_371, memorywre_371, 
        memoryro_362, memorywre_362, memoryro_363, memorywre_363, 
        memoryro_364, memorywre_364, memoryro_365, memorywre_365, 
        memoryro_366, memorywre_366, memoryro_357, memorywre_357, 
        memoryro_358, memorywre_358, memoryro_359, memorywre_359, 
        memoryro_360, memorywre_360, memoryro_361, memorywre_361, 
        memoryro_352, memorywre_352, memoryro_353, memorywre_353, 
        memoryro_354, memorywre_354, memoryro_355, memorywre_355, 
        memoryro_356, memorywre_356, memoryro_347, memorywre_347, 
        memoryro_348, memorywre_348, memoryro_349, memorywre_349, 
        memoryro_350, memorywre_350, memoryro_351, memorywre_351, 
        memoryro_342, memorywre_342, memoryro_343, memorywre_343, 
        memoryro_344, memorywre_344, memoryro_345, memorywre_345, 
        memoryro_346, memorywre_346, memoryro_337, memorywre_337, 
        memoryro_338, memorywre_338, memoryro_339, memorywre_339, 
        memoryro_340, memorywre_340, memoryro_341, memorywre_341, 
        memoryro_332, memorywre_332, memoryro_333, memorywre_333, 
        memoryro_334, memorywre_334, memoryro_335, memorywre_335, 
        memoryro_336, memorywre_336, memoryro_327, memorywre_327, 
        memoryro_328, memorywre_328, memoryro_329, memorywre_329, 
        memoryro_330, memorywre_330, memoryro_331, memorywre_331, 
        memoryro_322, memorywre_322, memoryro_323, memorywre_323, 
        memoryro_324, memorywre_324, memoryro_325, memorywre_325, 
        memoryro_326, memorywre_326, memoryro_317, memorywre_317, 
        memoryro_318, memorywre_318, memoryro_319, memorywre_319, 
        memoryro_320, memorywre_320, memoryro_321, memorywre_321, 
        memoryro_312, memorywre_312, memoryro_313, memorywre_313, 
        memoryro_314, memorywre_314, memoryro_315, memorywre_315, 
        memoryro_316, memorywre_316, memoryro_307, memorywre_307, 
        memoryro_308, memorywre_308, memoryro_309, memorywre_309, 
        memoryro_310, memorywre_310, memoryro_311, memorywre_311, 
        memoryro_302, memorywre_302, memoryro_303, memorywre_303, 
        memoryro_304, memorywre_304, memoryro_305, memorywre_305, 
        memoryro_306, memorywre_306, memoryro_297, memorywre_297, 
        memoryro_298, memorywre_298, memoryro_299, memorywre_299, 
        memoryro_300, memorywre_300, memoryro_301, memorywre_301, 
        memoryro_292, memorywre_292, memoryro_293, memorywre_293, 
        memoryro_294, memorywre_294, memoryro_295, memorywre_295, 
        memoryro_296, memorywre_296, memoryro_287, memorywre_287, 
        memoryro_288, memorywre_288, memoryro_289, memorywre_289, 
        memoryro_290, memorywre_290, memoryro_291, memorywre_291, 
        memoryro_282, memorywre_282, memoryro_283, memorywre_283, 
        memoryro_284, memorywre_284, memoryro_285, memorywre_285, 
        memoryro_286, memorywre_286, memoryro_277, memorywre_277, 
        memoryro_278, memorywre_278, memoryro_279, memorywre_279, 
        memoryro_280, memorywre_280, memoryro_281, memorywre_281, 
        memoryro_272, memorywre_272, memoryro_273, memorywre_273, 
        memoryro_274, memorywre_274, memoryro_275, memorywre_275, 
        memoryro_276, memorywre_276, memoryro_267, memorywre_267, 
        memoryro_268, memorywre_268, memoryro_269, memorywre_269, 
        memoryro_270, memorywre_270, memoryro_271, memorywre_271, 
        memoryro_262, memorywre_262, memoryro_263, memorywre_263, 
        memoryro_264, memorywre_264, memoryro_265, memorywre_265, 
        memoryro_266, memorywre_266, memoryro_257, memorywre_257, 
        memoryro_258, memorywre_258, memoryro_259, memorywre_259, 
        memoryro_260, memorywre_260, memoryro_261, memorywre_261, 
        memoryro_252, memorywre_252, memoryro_253, memorywre_253, 
        memoryro_254, memorywre_254, memoryro_255, memorywre_255, 
        memoryro_256, memorywre_256, memoryro_247, memorywre_247, 
        memoryro_248, memorywre_248, memoryro_249, memorywre_249, 
        memoryro_250, memorywre_250, memoryro_251, memorywre_251, 
        memoryro_242, memorywre_242, memoryro_243, memorywre_243, 
        memoryro_244, memorywre_244, memoryro_245, memorywre_245, 
        memoryro_246, memorywre_246, memoryro_237, memorywre_237, 
        memoryro_238, memorywre_238, memoryro_239, memorywre_239, 
        memoryro_240, memorywre_240, memoryro_241, memorywre_241, 
        memoryro_232, memorywre_232, memoryro_233, memorywre_233, 
        memoryro_234, memorywre_234, memoryro_235, memorywre_235, 
        memoryro_236, memorywre_236, memoryro_227, memorywre_227, 
        memoryro_228, memorywre_228, memoryro_229, memorywre_229, 
        memoryro_230, memorywre_230, memoryro_231, memorywre_231, 
        memoryro_222, memorywre_222, memoryro_223, memorywre_223, 
        memoryro_224, memorywre_224, memoryro_225, memorywre_225, 
        memoryro_226, memorywre_226, memoryro_217, memorywre_217, 
        memoryro_218, memorywre_218, memoryro_219, memorywre_219, 
        memoryro_220, memorywre_220, memoryro_221, memorywre_221, 
        memoryro_212, memorywre_212, memoryro_213, memorywre_213, 
        memoryro_214, memorywre_214, memoryro_215, memorywre_215, 
        memoryro_216, memorywre_216, memoryro_207, memorywre_207, 
        memoryro_208, memorywre_208, memoryro_209, memorywre_209, 
        memoryro_210, memorywre_210, memoryro_211, memorywre_211, 
        memoryro_202, memorywre_202, memoryro_203, memorywre_203, 
        memoryro_204, memorywre_204, memoryro_205, memorywre_205, 
        memoryro_206, memorywre_206, memoryro_197, memorywre_197, 
        memoryro_198, memorywre_198, memoryro_199, memorywre_199, 
        memoryro_200, memorywre_200, memoryro_201, memorywre_201, 
        memoryro_192, memorywre_192, memoryro_193, memorywre_193, 
        memoryro_194, memorywre_194, memoryro_195, memorywre_195, 
        memoryro_196, memorywre_196, memoryro_187, memorywre_187, 
        memoryro_188, memorywre_188, memoryro_189, memorywre_189, 
        memoryro_190, memorywre_190, memoryro_191, memorywre_191, 
        memoryro_182, memorywre_182, memoryro_183, memorywre_183, 
        memoryro_184, memorywre_184, memoryro_185, memorywre_185, 
        memoryro_186, memorywre_186, memoryro_177, memorywre_177, 
        memoryro_178, memorywre_178, memoryro_179, memorywre_179, 
        memoryro_180, memorywre_180, memoryro_181, memorywre_181, 
        memoryro_172, memorywre_172, memoryro_173, memorywre_173, 
        memoryro_174, memorywre_174, memoryro_175, memorywre_175, 
        memoryro_176, memorywre_176, memoryro_167, memorywre_167, 
        memoryro_168, memorywre_168, memoryro_169, memorywre_169, 
        memoryro_170, memorywre_170, memoryro_171, memorywre_171, 
        memoryro_162, memorywre_162, memoryro_163, memorywre_163, 
        memoryro_164, memorywre_164, memoryro_165, memorywre_165, 
        memoryro_166, memorywre_166, memoryro_157, memorywre_157, 
        memoryro_158, memorywre_158, memoryro_159, memorywre_159, 
        memoryro_160, memorywre_160, memoryro_161, memorywre_161, 
        memoryro_152, memorywre_152, memoryro_153, memorywre_153, 
        memoryro_154, memorywre_154, memoryro_155, memorywre_155, 
        memoryro_156, memorywre_156, memoryro_147, memorywre_147, 
        memoryro_148, memorywre_148, memoryro_149, memorywre_149, 
        memoryro_150, memorywre_150, memoryro_151, memorywre_151, 
        memoryro_142, memorywre_142, memoryro_143, memorywre_143, 
        memoryro_144, memorywre_144, memoryro_145, memorywre_145, 
        memoryro_146, memorywre_146, memoryro_137, memorywre_137, 
        memoryro_138, memorywre_138, memoryro_139, memorywre_139, 
        memoryro_140, memorywre_140, memoryro_141, memorywre_141, 
        memoryro_132, memorywre_132, memoryro_133, memorywre_133, 
        memoryro_134, memorywre_134, memoryro_135, memorywre_135, 
        memoryro_136, memorywre_136, memoryro_127, memorywre_127, 
        memoryro_128, memorywre_128, memoryro_129, memorywre_129, 
        memoryro_130, memorywre_130, memoryro_131, memorywre_131, 
        memoryro_122, memorywre_122, memoryro_123, memorywre_123, 
        memoryro_124, memorywre_124, memoryro_125, memorywre_125, 
        memoryro_126, memorywre_126, memoryro_117, memorywre_117, 
        memoryro_118, memorywre_118, memoryro_119, memorywre_119, 
        memoryro_120, memorywre_120, memoryro_121, memorywre_121, 
        memoryro_112, memorywre_112, memoryro_113, memorywre_113, 
        memoryro_114, memorywre_114, memoryro_115, memorywre_115, 
        memoryro_116, memorywre_116, memoryro_107, memorywre_107, 
        memoryro_108, memorywre_108, memoryro_109, memorywre_109, 
        memoryro_110, memorywre_110, memoryro_111, memorywre_111, 
        memoryro_102, memorywre_102, memoryro_103, memorywre_103, 
        memoryro_104, memorywre_104, memoryro_105, memorywre_105, 
        memoryro_106, memorywre_106, memoryro_97, memorywre_97, 
        memoryro_98, memorywre_98, memoryro_99, memorywre_99, 
        memoryro_100, memorywre_100, memoryro_101, memorywre_101, 
        memoryro_92, memorywre_92, memoryro_93, memorywre_93, 
        memoryro_94, memorywre_94, memoryro_95, memorywre_95, 
        memoryro_96, memorywre_96, memoryro_87, memorywre_87, 
        memoryro_88, memorywre_88, memoryro_89, memorywre_89, 
        memoryro_90, memorywre_90, memoryro_91, memorywre_91, 
        memoryro_82, memorywre_82, memoryro_83, memorywre_83, 
        memoryro_84, memorywre_84, memoryro_85, memorywre_85, 
        memoryro_86, memorywre_86, memoryro_77, memorywre_77, 
        memoryro_78, memorywre_78, memoryro_79, memorywre_79, 
        memoryro_80, memorywre_80, memoryro_81, memorywre_81, 
        memoryro_72, memorywre_72, memoryro_73, memorywre_73, 
        memoryro_74, memorywre_74, memoryro_75, memorywre_75, 
        memoryro_76, memorywre_76, memoryro_67, memorywre_67, 
        memoryro_68, memorywre_68, memoryro_69, memorywre_69, 
        memoryro_70, memorywre_70, memoryro_71, memorywre_71, 
        memoryro_62, memorywre_62, memoryro_63, memorywre_63, 
        memoryro_64, memorywre_64, memoryro_65, memorywre_65, 
        memoryro_66, memorywre_66, memoryro_57, memorywre_57, 
        memoryro_58, memorywre_58, memoryro_59, memorywre_59, 
        memoryro_60, memorywre_60, memoryro_61, memorywre_61, 
        memoryro_52, memorywre_52, memoryro_53, memorywre_53, 
        memoryro_54, memorywre_54, memoryro_55, memorywre_55, 
        memoryro_56, memorywre_56, memoryro_47, memorywre_47, 
        memoryro_48, memorywre_48, memoryro_49, memorywre_49, 
        memoryro_50, memorywre_50, memoryro_51, memorywre_51, 
        memoryro_42, memorywre_42, memoryro_43, memorywre_43, 
        memoryro_44, memorywre_44, memoryro_45, memorywre_45, 
        memoryro_46, memorywre_46, memoryro_37, memorywre_37, 
        memoryro_38, memorywre_38, memoryro_39, memorywre_39, 
        memoryro_40, memorywre_40, memoryro_41, memorywre_41, 
        memoryro_32, memorywre_32, memoryro_33, memorywre_33, 
        memoryro_34, memorywre_34, memoryro_35, memorywre_35, 
        memoryro_36, memorywre_36, memoryro_27, memorywre_27, 
        memoryro_28, memorywre_28, memoryro_29, memorywre_29, 
        memoryro_30, memorywre_30, memoryro_31, memorywre_31, 
        memoryro_22, memorywre_22, memoryro_23, memorywre_23, 
        memoryro_24, memorywre_24, memoryro_25, memorywre_25, 
        memoryro_26, memorywre_26, memoryro_17, memorywre_17, 
        memoryro_18, memorywre_18, memoryro_19, memorywre_19, 
        memoryro_20, memorywre_20, memoryro_21, memorywre_21, 
        memoryro_12, memorywre_12, memoryro_13, memorywre_13, 
        memoryro_14, memorywre_14, memoryro_15, memorywre_15, 
        memoryro_16, memorywre_16, memoryro_7, memorywre_7, 
        memoryro_8, memorywre_8, memoryro_9, memorywre_9, 
        memoryro_10, memorywre_10, memoryro_11, memorywre_11, 
        memoryro_2, memorywre_2, memoryro_3, memorywre_3, 
        memoryro_4, memorywre_4, memoryro_5, memorywre_5, 
        memoryro_6, memorywre_6, memoryro_0, memorywre_0, 
        memoryro_1, memorywre_1, memory_memory_0_0_en_Z, 
        dout_1_sqmuxa_Z, memory_memory_0_0_sr_Z, memoryror_i, 
        memorya116_1_Z, memorya20_0_Z, memorya20_6_Z, 
        memorya36_1_Z, memorya36_6_Z, memorya102_1_Z, 
        memorya16_0_Z, memorya117_1_Z, memorya5_0_Z, memorya4_6_Z, 
        memorya21_0_Z, memorya57_3_Z, memorya9_0_Z, memorya8_0_Z, 
        memorya368_6_Z, memorya368_0_Z, memorya305_2_Z, 
        memorya298_6_Z, memorya266_0_Z, memorya499_5_Z, 
        memorya435_6_Z, memorya193_2_Z, memorya369_5_Z, 
        memorya3_0_Z, memorya68_3_Z, memorya273_4_Z, 
        memorya128_0_Z, memorya403_2_Z, memorya273_6_Z, 
        memorya432_0_Z, memorya162_2_Z, memorya264_6_Z, 
        memorya42_0_Z, memorya395_2_Z, memorya227_0_Z, 
        memorya101_5_Z, memorya464_0_Z, memorya441_6_Z, 
        memorya264_1_Z, memorya268_6_Z, memorya261_0_Z, 
        memorya292_6_Z, memorya211_3_Z, memorya331_5_Z, 
        memorya199_0_Z, memorya455_5_Z, memorya167_3_Z, 
        memorya102_5_Z, memorya463_5_Z, memorya111_0_Z, 
        memorya102_4_Z, memorya124_0_Z, memorya380_5_Z, 
        memorya84_2_Z, memorya52_2_Z, memorya45_6_Z, 
        memorya12_0_Z, memorya68_2_Z, memorya121_4_Z, 
        memorya315_5_Z, memorya362_1_Z, memorya10_0_Z, 
        memorya116_4_Z, memorya503_5_Z, memorya379_1_Z, 
        memorya35_0_Z, memorya354_1_Z, memorya370_1_Z, 
        memorya86_2_Z, memorya83_6_Z, memorya54_2_Z, 
        memorya51_6_Z, memorya372_6_Z, memorya482_2_Z, 
        memorya468_Z, memorya340_6_Z, memorya212_Z, 
        memorya320_6_Z, memorya498_3_Z, memorya384_Z, 
        memorya444_Z, memorya434_2_Z, memorya436_Z, memorya93_0, 
        memorya117_Z, memorya245_Z, memorya211_0_Z, memorya213_Z, 
        memorya125_2_Z, memorya376_6_Z, memorya440_Z, 
        memorya345_6_Z, memorya121_1_Z, memorya345_Z, 
        memorya473_Z, memorya498_6_Z, memorya474_Z, memorya68_4_Z, 
        memorya90_Z, memorya364_1_Z, memorya204_6_Z, memorya204_Z, 
        memorya364_6_Z, memorya460_Z, memorya428_Z, memorya93_Z, 
        memorya116_2_Z, memorya125_Z, memorya253_Z, 
        memorya368_4_Z, memorya96_Z, memorya353_1_Z, 
        memorya353_6_Z, memorya225_Z, memorya447_Z, memorya479_Z, 
        memorya383_Z, memorya503_Z, memorya507_Z, memorya495_Z, 
        memorya126_5_Z, memorya510_Z, memorya381_5_Z, 
        memorya509_Z, memorya480_Z, memorya504_6_Z, memorya476_Z, 
        memorya92_Z, memorya250_Z, memorya442_Z, memorya52_4, 
        memorya58_Z, memorya289_4_Z, memorya160_Z, memorya128, 
        memorya391_2_Z, memorya132_Z, memorya386_1_Z, 
        memorya130_Z, memorya369_3_Z, memorya261_Z, memorya256_Z, 
        memorya369_Z, memorya481_5_Z, memorya481_Z, 
        memorya304_4_Z, memorya63_0, memorya176_Z, memorya77_2_Z, 
        memorya206_Z, memorya333_6_Z, memorya333_Z, memorya205_Z, 
        memorya45_2_Z, memorya45_Z, memorya109_Z, memorya236_0_Z, 
        memorya237_Z, memorya121_Z, memorya441_Z, memorya342_6_Z, 
        memorya342_Z, memorya214_Z, memorya68_1_Z, memorya68_Z, 
        memorya66_1_Z, memorya66_Z, memorya71_Z, memorya4_3_Z, 
        memoryror_483, memoryror_504_1, memoryror_482, 
        memoryror_481, memoryror_504, memoryror_387, 
        memoryror_386, memoryror_385, memoryror_384, memorya4_0_Z, 
        memorya13_0_Z, memorya2_0_Z, memorya1_0_Z, memorya11_0_Z, 
        memorya7_0_Z, memorya19_0_Z, memorya258_0_Z, 
        memorya257_0_Z, memorya31_0_Z, memorya223_0_Z, 
        memorya79_0_Z, memorya47_0_Z, memorya126_0_Z, 
        memorya55_0_Z, memorya67_2_Z, memorya193_1_Z, 
        memorya385_1_Z, memorya415_4_Z, memorya463_4_Z, 
        memorya487_4_Z, memorya318_4_Z, memorya316_4_Z, 
        memorya379_4_Z, memorya312_4_Z, memorya278_2_Z, 
        memorya260_1_Z, memorya370_3_Z, memorya354_3_Z, 
        memorya369_1_Z, memorya368_2_Z, memorya46_3_Z, 
        memorya30_3_Z, memorya45_3_Z, memorya29_3_Z, 
        memorya41_3_Z, memorya25_3_Z, memorya117_3_Z, 
        memorya37_2_Z, memorya102_3_Z, memorya84_3_Z, 
        memorya20_3_Z, memorya87_0, memorya143_0_Z, memorya56_0_Z, 
        memorya52_0_Z, memorya233_0_Z, memorya280_0_Z, 
        memorya276_0_Z, memorya268_0_Z, memorya361_6_Z, 
        memorya156_5_Z, memorya100_6_Z, memorya339_6_Z, 
        memorya355_6_Z, memorya436_5_Z, memorya197_6_Z, 
        memorya118_5_Z, memorya373_5_Z, memorya421_6_Z, 
        memorya213_5_Z, memorya149_5_Z, memorya336_6_Z, 
        memorya326_6_Z, memorya440_5_Z, memorya393_6_Z, 
        memorya345_5_Z, memorya474_5_Z, memorya154_5_Z, 
        memorya202_6_Z, memorya428_5_Z, memorya142_5_Z, 
        memorya98_6_Z, memorya395_5_Z, memorya487_5_Z, 
        memorya391_6_Z, memorya270_6_Z, memorya348_5_Z, 
        memorya299_5_Z, memorya378_5_Z, memorya362_6_Z, 
        memorya344_6_Z, memorya296_6_Z, memorya280_6_Z, 
        memorya360_6_Z, memorya294_6_Z, memorya278_6_Z, 
        memorya358_6_Z, memorya356_6_Z, memorya370_6_Z, 
        memorya338_6_Z, memorya306_6_Z, memorya354_6_Z, 
        memorya289_6_Z, memorya257_6_Z, memorya369_6_Z, 
        memorya304_6_Z, memorya78_5_Z, memorya110_5_Z, 
        memorya77_5_Z, memorya45_5_Z, memorya105_6_Z, 
        memorya121_5_Z, memorya86_5_Z, memorya68_6_Z, memorya4_Z, 
        memorya20, memorya36, memorya52_Z, memorya84_Z, 
        memorya116_Z, memorya6_Z, memorya22, memorya38_Z, 
        memorya54_Z, memorya86_Z, memorya102_Z, memorya70_Z, 
        memorya5, memorya21, memorya37_Z, memorya53_Z, 
        memorya85_Z, memorya101_Z, memorya69_Z, memorya9, 
        memorya25_Z, memorya41_Z, memorya57_Z, memorya89_Z, 
        memorya105_Z, memorya73_Z, memorya13_Z, memorya29_Z, 
        memorya61_Z, memorya77_Z, memorya14, memorya30_Z, 
        memorya46_Z, memorya62_Z, memorya94_Z, memorya110_Z, 
        memorya78_Z, memorya304_Z, memorya320_Z, memorya368, 
        memorya257_Z, memorya273_Z, memorya289_Z, memorya305_Z, 
        memorya337_Z, memorya353_Z, memorya354_Z, memorya258_Z, 
        memorya274_Z, memorya290_Z, memorya306_Z, memorya338_Z, 
        memorya370_Z, memorya356_Z, memorya260_Z, memorya276_Z, 
        memorya292_Z, memorya308_Z, memorya340_Z, memorya372_Z, 
        memorya358_Z, memorya262_Z, memorya278_Z, memorya294_Z, 
        memorya310_Z, memorya374_Z, memorya264_Z, memorya280_Z, 
        memorya296_Z, memorya312_Z, memorya344_Z, memorya360_Z, 
        memorya376_Z, memorya362_Z, memorya266_Z, memorya282_Z, 
        memorya298, memorya314_Z, memorya346_Z, memorya378_Z, 
        memorya267_Z, memorya299_Z, memorya315_Z, memorya331_Z, 
        memorya347_Z, memorya363_Z, memorya364_Z, memorya268_Z, 
        memorya284_Z, memorya300_Z, memorya316_Z, memorya348_Z, 
        memorya380_Z, memorya366_Z, memorya270_Z, memorya286_Z, 
        memorya302_Z, memorya318_Z, memorya350_Z, memorya382_Z, 
        memorya386_Z, memorya402_Z, memorya418_Z, memorya434_Z, 
        memorya466_Z, memorya482_Z, memorya498_Z, memorya387_Z, 
        memorya403_Z, memorya419_Z, memorya435, memorya451_Z, 
        memorya467_Z, memorya483_Z, memorya499_Z, memorya455_Z, 
        memorya391_Z, memorya407_Z, memorya423_Z, memorya471_Z, 
        memorya487_Z, memorya395_Z, memorya411_Z, memorya427_Z, 
        memorya459_Z, memorya491_Z, memorya475_Z, memorya463_Z, 
        memorya399_Z, memorya415_Z, memorya431_Z, memorya385_Z, 
        memorya433_Z, memorya465_Z, memorya193_Z, memorya321_Z, 
        memorya129_Z, memorya145_Z, memorya161_Z, memorya177_Z, 
        memorya209_Z, memorya241, memorya162_Z, memorya98_Z, 
        memorya97_Z, memorya65_Z, memorya194_Z, memorya226_Z, 
        memorya242_Z, memorya450_Z, memorya144, memorya432, 
        memorya400_Z, memorya351_Z, memorya64_Z, memorya352_Z, 
        memorya334_Z, memorya142_Z, memorya158_Z, memorya190_Z, 
        memorya446_Z, memorya141_Z, memorya173_Z, memorya189_Z, 
        memorya221_Z, memorya429_Z, memorya430_Z, memorya349_Z, 
        memorya174_Z, memorya126_Z, memorya188_Z, memorya220_Z, 
        memorya252_Z, memorya202_Z, memorya234_Z, memorya138, 
        memorya154_Z, memorya186_Z, memorya218_Z, memorya330_Z, 
        memorya137, memorya153_Z, memorya169_Z, memorya185_Z, 
        memorya217_Z, memorya425_Z, memorya424_Z, memorya377_Z, 
        memorya170_Z, memorya106_Z, memorya74_Z, memorya393_Z, 
        memorya409_Z, memorya328_Z, memorya136, memorya152_Z, 
        memorya184_Z, memorya408_Z, memorya392_Z, memorya343_Z, 
        memorya168_Z, memorya104_Z, memorya72_Z, memorya166_Z, 
        memorya326_Z, memorya134_Z, memorya150_Z, memorya182_Z, 
        memorya438_Z, memorya336_Z, memorya416_Z, memorya133_Z, 
        memorya149_Z, memorya165_Z, memorya181_Z, memorya421_Z, 
        memorya437_Z, memorya422_Z, memorya373_Z, memorya341_Z, 
        memorya118_Z, memorya197_Z, memorya229, memorya420_Z, 
        memorya324_Z, memorya148_Z, memorya164_Z, memorya228_Z, 
        memorya259_Z, memorya275_Z, memorya307_Z, memorya323_Z, 
        memorya339_Z, memorya355_Z, memorya371_Z, memorya131_Z, 
        memorya147_Z, memorya163_Z, memorya179_Z, memorya211_Z, 
        memorya243_Z, memorya404_Z, memorya388_Z, memorya180_Z, 
        memorya100_Z, memorya67_Z, memorya99_Z, memorya227_Z, 
        memorya291_Z, memorya359_Z, memorya327_Z, memorya183_Z, 
        memorya167_Z, memorya135_Z, memorya219_Z, memorya187_Z, 
        memorya171_Z, memorya139_Z, memorya236_Z, memorya172_Z, 
        memorya156_Z, memorya140_Z, memorya367_Z, memorya335_Z, 
        memorya191_Z, memorya175_Z, memorya159_Z, memorya143_Z, 
        memorya210_Z, memorya178_Z, memorya146_Z, memorya494_Z, 
        memorya478_Z, memorya462_Z, memorya493_Z, memorya477_Z, 
        memorya461_Z, memorya508_Z, memorya492_Z, memorya505_Z, 
        memorya489_Z, memorya457_Z, memorya504_Z, memorya488_Z, 
        memorya472_Z, memorya456_Z, memorya502_Z, memorya486_Z, 
        memorya470_Z, memorya454_Z, memorya501_Z, memorya485_Z, 
        memorya469_Z, memorya453_Z, memorya500_Z, memorya484_Z, 
        memorya452_Z, memorya496_Z, memorya464, memorya448_Z, 
        memorya414_Z, memorya398_Z, memorya413_Z, memorya397_Z, 
        memorya412_Z, memorya396_Z, memorya506_Z, memorya490_Z, 
        memorya458_Z, memorya426_Z, memorya410_Z, memorya394_Z, 
        memorya406_Z, memorya390_Z, memorya405_Z, memorya389_Z, 
        memorya497, memorya449_Z, memorya417_Z, memorya401_Z, 
        memorya319_Z, memorya303_Z, memorya287_Z, memorya271_Z, 
        memorya365_Z, memorya317_Z, memorya301_Z, memorya269, 
        memorya332_Z, memorya361_Z, memorya329_Z, memorya313_Z, 
        memorya297_Z, memorya281_Z, memorya265_Z, memorya311_Z, 
        memorya295_Z, memorya263_Z, memorya357_Z, memorya325_Z, 
        memorya309_Z, memorya293, memorya277_Z, memorya322_Z, 
        memorya288_Z, memorya272_Z, memorya239_Z, memorya223_Z, 
        memorya207_Z, memorya254_Z, memorya238_Z, memorya222_Z, 
        memorya235_Z, memorya203, memorya249_Z, memorya233_Z, 
        memorya201_Z, memorya248_Z, memorya232_Z, memorya216_Z, 
        memorya200_Z, memorya231_Z, memorya215_Z, memorya199, 
        memorya246_Z, memorya230, memorya198_Z, memorya244_Z, 
        memorya196_Z, memorya208_Z, memorya111, memorya79_Z, 
        memorya108_Z, memorya76_Z, memorya107_Z, memorya75_Z, 
        memorya103_Z, memorya127_Z, memorya95_Z, memorya63_Z, 
        memorya47_Z, memorya31_Z, memorya15, memorya124, 
        memorya60_Z, memorya44, memorya28_Z, memorya12, 
        memorya123, memorya91_Z, memorya59_Z, memorya43_Z, 
        memorya27_Z, memorya11_Z, memorya122_Z, memorya42_Z, 
        memorya26_Z, memorya10, memorya120_Z, memorya88_Z, 
        memorya56_Z, memorya40_Z, memorya24_Z, memorya8, 
        memorya119, memorya87_Z, memorya55_Z, memorya39_Z, 
        memorya23_Z, memorya7_Z, memorya115_Z, memorya83_Z, 
        memorya51_Z, memorya35, memorya19_Z, memorya3, 
        memorya114_Z, memorya82_Z, memorya50_Z, memorya34, 
        memorya18, memorya2_Z, memorya113_Z, memorya81_Z, 
        memorya49_Z, memorya33_Z, memorya17_Z, memorya1_Z, 
        memorya112_Z, memorya80, memorya48, memorya32_Z, 
        memorya16, memorya0, memorya192_Z, memorya224_Z, 
        memorya240_Z, memorya247, memorya279_Z, memorya285_Z, 
        memorya155_Z, memorya251, memorya151_Z, memorya195_Z, 
        memorya375_Z, memorya381_Z, memorya445_Z, memorya157_Z, 
        memorya443_Z, memorya439_Z, memorya379_Z, memorya283_Z, 
        memorya255_Z, memorya511_Z, memoryror_255, memoryror_254, 
        memoryror_253, memoryror_252, memoryror_251, 
        memoryror_250, memoryror_249, memoryror_248, 
        memoryror_247, memoryror_246, memoryror_245, 
        memoryror_244, memoryror_243, memoryror_242, 
        memoryror_241, memoryror_240, memoryror_239, 
        memoryror_238, memoryror_237, memoryror_236, 
        memoryror_235, memoryror_234, memoryror_233, 
        memoryror_232, memoryror_231, memoryror_230, 
        memoryror_229, memoryror_228, memoryror_227, 
        memoryror_226, memoryror_225, memoryror_224, 
        memoryror_223, memoryror_222, memoryror_221, 
        memoryror_220, memoryror_219, memoryror_218, 
        memoryror_217, memoryror_216, memoryror_215, 
        memoryror_214, memoryror_213, memoryror_212, 
        memoryror_211, memoryror_210, memoryror_209, 
        memoryror_208, memoryror_207, memoryror_206, 
        memoryror_205, memoryror_204, memoryror_203, 
        memoryror_202, memoryror_201, memoryror_200, 
        memoryror_199, memoryror_198, memoryror_197, 
        memoryror_196, memoryror_195, memoryror_194, 
        memoryror_193, memoryror_192, memoryror_191, 
        memoryror_190, memoryror_189, memoryror_188, 
        memoryror_187, memoryror_186, memoryror_185, 
        memoryror_184, memoryror_183, memoryror_182, 
        memoryror_181, memoryror_180, memoryror_179, 
        memoryror_178, memoryror_177, memoryror_176, 
        memoryror_175, memoryror_174, memoryror_173, 
        memoryror_172, memoryror_171, memoryror_170, 
        memoryror_169, memoryror_168, memoryror_167, 
        memoryror_166, memoryror_165, memoryror_164, 
        memoryror_163, memoryror_162, memoryror_161, 
        memoryror_160, memoryror_159, memoryror_158, 
        memoryror_157, memoryror_156, memoryror_155, 
        memoryror_154, memoryror_153, memoryror_152, 
        memoryror_151, memoryror_150, memoryror_149, 
        memoryror_148, memoryror_147, memoryror_146, 
        memoryror_145, memoryror_144, memoryror_143, 
        memoryror_142, memoryror_141, memoryror_140, 
        memoryror_139, memoryror_138, memoryror_137, 
        memoryror_136, memoryror_135, memoryror_134, 
        memoryror_133, memoryror_132, memoryror_131, 
        memoryror_130, memoryror_129, memoryror_128, 
        memoryror_127, memoryror_126, memoryror_125, 
        memoryror_124, memoryror_123, memoryror_122, 
        memoryror_121, memoryror_120, memoryror_119, 
        memoryror_118, memoryror_117, memoryror_116, 
        memoryror_115, memoryror_114, memoryror_113, 
        memoryror_112, memoryror_111, memoryror_110, 
        memoryror_109, memoryror_108, memoryror_107, 
        memoryror_106, memoryror_105, memoryror_104, 
        memoryror_103, memoryror_102, memoryror_101, 
        memoryror_100, memoryror_99, memoryror_98, memoryror_97, 
        memoryror_96, memoryror_95, memoryror_94, memoryror_93, 
        memoryror_92, memoryror_91, memoryror_90, memoryror_89, 
        memoryror_88, memoryror_87, memoryror_86, memoryror_85, 
        memoryror_84, memoryror_83, memoryror_82, memoryror_81, 
        memoryror_80, memoryror_79, memoryror_78, memoryror_77, 
        memoryror_76, memoryror_75, memoryror_74, memoryror_73, 
        memoryror_72, memoryror_71, memoryror_70, memoryror_69, 
        memoryror_68, memoryror_67, memoryror_66, memoryror_65, 
        memoryror_64, memoryror_63, memoryror_62, memoryror_61, 
        memoryror_60, memoryror_59, memoryror_58, memoryror_57, 
        memoryror_56, memoryror_55, memoryror_54, memoryror_53, 
        memoryror_52, memoryror_51, memoryror_50, memoryror_49, 
        memoryror_48, memoryror_47, memoryror_46, memoryror_45, 
        memoryror_44, memoryror_43, memoryror_42, memoryror_41, 
        memoryror_40, memoryror_39, memoryror_38, memoryror_37, 
        memoryror_36, memoryror_35, memoryror_34, memoryror_33, 
        memoryror_32, memoryror_31, memoryror_30, memoryror_29, 
        memoryror_28, memoryror_27, memoryror_26, memoryror_25, 
        memoryror_24, memoryror_23, memoryror_22, memoryror_21, 
        memoryror_20, memoryror_19, memoryror_18, memoryror_17, 
        memoryror_16, memoryror_15, memoryror_14, memoryror_13, 
        memoryror_12, memoryror_11, memoryror_10, memoryror_9, 
        memoryror_8, memoryror_7, memoryror_6, memoryror_5, 
        memoryror_4, memoryror_3, memoryror_2, memoryror_1, 
        memoryror_0, memoryror_447, memoryror_446, memoryror_445, 
        memoryror_444, memoryror_443, memoryror_442, 
        memoryror_441, memoryror_440, memoryror_439, 
        memoryror_438, memoryror_437, memoryror_436, 
        memoryror_435, memoryror_434, memoryror_433, 
        memoryror_432, memoryror_431, memoryror_430, 
        memoryror_429, memoryror_428, memoryror_427, 
        memoryror_426, memoryror_425, memoryror_424, 
        memoryror_423, memoryror_422, memoryror_421, 
        memoryror_420, memoryror_419, memoryror_418, 
        memoryror_417, memoryror_416, memoryror_415, 
        memoryror_414, memoryror_413, memoryror_412, 
        memoryror_411, memoryror_410, memoryror_409, 
        memoryror_408, memoryror_407, memoryror_406, 
        memoryror_405, memoryror_404, memoryror_403, 
        memoryror_402, memoryror_401, memoryror_400, 
        memoryror_399, memoryror_398, memoryror_397, 
        memoryror_396, memoryror_395, memoryror_394, 
        memoryror_393, memoryror_392, memoryror_391, 
        memoryror_390, memoryror_389, memoryror_388, 
        memoryror_495, memoryror_494, memoryror_493, 
        memoryror_492, memoryror_491, memoryror_490, 
        memoryror_489, memoryror_488, memoryror_487, 
        memoryror_486, memoryror_485, memoryror_484, 
        memoryror_507, memoryror_506, memoryror_505, NC0
         : std_logic;

begin 

    InternalDataFromMem(31) <= \InternalDataFromMem\(31);
    InternalDataFromMem(30) <= \InternalDataFromMem\(30);
    InternalDataFromMem(29) <= \InternalDataFromMem\(29);
    InternalDataFromMem(28) <= \InternalDataFromMem\(28);
    InternalDataFromMem(27) <= \InternalDataFromMem\(27);
    InternalDataFromMem(26) <= \InternalDataFromMem\(26);
    InternalDataFromMem(25) <= \InternalDataFromMem\(25);
    InternalDataFromMem(24) <= \InternalDataFromMem\(24);
    InternalDataFromMem(23) <= \InternalDataFromMem\(23);
    InternalDataFromMem(22) <= \InternalDataFromMem\(22);
    InternalDataFromMem(21) <= \InternalDataFromMem\(21);
    InternalDataFromMem(20) <= \InternalDataFromMem\(20);
    InternalDataFromMem(19) <= \InternalDataFromMem\(19);
    InternalDataFromMem(18) <= \InternalDataFromMem\(18);
    InternalDataFromMem(17) <= \InternalDataFromMem\(17);
    InternalDataFromMem(16) <= \InternalDataFromMem\(16);
    InternalDataFromMem(15) <= \InternalDataFromMem\(15);
    InternalDataFromMem(14) <= \InternalDataFromMem\(14);
    InternalDataFromMem(13) <= \InternalDataFromMem\(13);
    InternalDataFromMem(12) <= \InternalDataFromMem\(12);
    InternalDataFromMem(11) <= \InternalDataFromMem\(11);
    InternalDataFromMem(10) <= \InternalDataFromMem\(10);
    InternalDataFromMem(9) <= \InternalDataFromMem\(9);
    InternalDataFromMem(8) <= \InternalDataFromMem\(8);
    InternalDataFromMem(7) <= \InternalDataFromMem\(7);
    InternalDataFromMem(6) <= \InternalDataFromMem\(6);
    InternalDataFromMem(5) <= \InternalDataFromMem\(5);
    InternalDataFromMem(4) <= \InternalDataFromMem\(4);
    InternalDataFromMem(3) <= \InternalDataFromMem\(3);
    InternalDataFromMem(2) <= \InternalDataFromMem\(2);
    InternalDataFromMem(1) <= \InternalDataFromMem\(1);
    InternalDataFromMem(0) <= \InternalDataFromMem\(0);

    memory_memory_0_0_sr_RNO_52 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_94, B => memoryror_95, C => 
        memoryror_92, D => memoryror_93, Y => memoryror_407);
    
    memory_memory_0_0_sr_RNO_47 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_130, B => memoryror_131, C => 
        memoryror_129, D => memoryror_128, Y => memoryror_416);
    
    memorya109_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya117_3_Z, B => InternalAddr2Memory(8), 
        Y => memorya93_0);
    
    memoryrff_48 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_48, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_48);
    
    memorya173 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya193_2_Z, B => memorya45_5_Z, C => 
        InternalAddr2Memory(8), D => memorya289_4_Z, Y => 
        memorya173_Z);
    
    memorya386 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya370_3_Z, B => memorya320_6_Z, C => 
        InternalAddr2Memory(6), D => memorya386_1_Z, Y => 
        memorya386_Z);
    
    memorya60 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya380_5_Z, B => memorya20_0_Z, C => 
        memorya52_4, Y => memorya60_Z);
    
    memorya78 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya46_3_Z, C
         => memorya68_4_Z, D => memorya78_5_Z, Y => memorya78_Z);
    
    memoryrff_262 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_262, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_262);
    
    memoryrff_72 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_72, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_72);
    
    memory_memory_0_0_sr_RNO_262 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_28, B => memoryro_508, C => 
        memorya508_Z, D => memorya28_Z, Y => memoryror_116);
    
    \memory_memory_0_0_OLDA[22]\ : SLE
      port map(D => \InternalDataFromMem\(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(22));
    
    memoryrff_285 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_285, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_285);
    
    memoryrff_68_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya68_Z, B => WriteEnable, Y => 
        memorywre_68);
    
    memoryrff_408_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya408_Z, B => WriteEnable, Y => 
        memorywre_408);
    
    memoryrff_20 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_20, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_20);
    
    memorya156_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya403_2_Z, B => memorya364_1_Z, Y => 
        memorya156_5_Z);
    
    \memory_memory_0_0_OLDA[16]\ : SLE
      port map(D => \InternalDataFromMem\(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(16));
    
    memoryrff_459 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_459, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_459);
    
    memoryrff_260_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya260_Z, B => WriteEnable, Y => 
        memorywre_260);
    
    memoryrff_204 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_204, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_204);
    
    memorya285 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya273_4_Z, 
        C => memorya369_3_Z, D => memorya381_5_Z, Y => 
        memorya285_Z);
    
    memory_memory_0_0_sr_RNO_144 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_243, B => memoryro_371, C => 
        memorya371_Z, D => memorya243_Z, Y => memoryror_248);
    
    memorya403 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_1_Z, B => InternalAddr2Memory(6), 
        C => memorya339_6_Z, D => memorya403_2_Z, Y => 
        memorya403_Z);
    
    memorya102 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya102_3_Z, 
        C => memorya102_4_Z, D => memorya102_5_Z, Y => 
        memorya102_Z);
    
    memory_memory_0_0_sr_RNO_82 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_31, B => memoryror_29, C => 
        memoryror_30, D => memoryror_28, Y => memoryror_391);
    
    memoryrff_479 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_479, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_479);
    
    memoryrff_223 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_223, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_223);
    
    memory_memory_0_0_sr_RNO_323 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_294, B => memoryro_38, C => 
        memorya294_Z, D => memorya38_Z, Y => memoryror_42);
    
    memoryrff_95_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya95_Z, B => WriteEnable, Y => 
        memorywre_95);
    
    memoryrff_35_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya379_1_Z, B => WriteEnable, C => 
        memorya36_6_Z, D => memorya35_0_Z, Y => memorywre_35);
    
    memoryrff_201_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya201_Z, B => WriteEnable, Y => 
        memorywre_201);
    
    memoryrff_67_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya67_Z, B => WriteEnable, Y => 
        memorywre_67);
    
    memory_memory_0_0_sr_RNO_101 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_98, B => memoryro_290, C => 
        memorya290_Z, D => memorya98_Z, Y => memoryror_224);
    
    memorya503_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya379_1_Z, B => memorya116_1_Z, Y => 
        memorya503_5_Z);
    
    memorya292_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya289_4_Z, B => memorya84_3_Z, Y => 
        memorya292_6_Z);
    
    memoryrff_3_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya379_1_Z, B => WriteEnable, C => 
        memorya4_6_Z, D => memorya3_0_Z, Y => memorywre_3);
    
    memorya354_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(1), Y => memorya354_1_Z);
    
    memoryrff_413_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya413_Z, B => WriteEnable, Y => 
        memorywre_413);
    
    memoryrff_111 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_111, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_111);
    
    memory_memory_0_0_sr_RNO_189 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_248, B => memoryro_264, C => 
        memorya264_Z, D => memorya248_Z, Y => memoryror_143);
    
    memorya79_0 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(4), Y => memorya79_0_Z);
    
    memory_memory_0_0_sr_RNO_180 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_324, B => memoryro_132, C => 
        memorya324_Z, D => memorya132_Z, Y => memoryror_137);
    
    memorya125_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(3), Y => memorya125_2_Z);
    
    memoryrff_303_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya303_Z, B => WriteEnable, Y => 
        memorywre_303);
    
    memorya183 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya304_4_Z, 
        C => memorya434_2_Z, D => memorya503_5_Z, Y => 
        memorya183_Z);
    
    memorya368_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(6), Y => memorya368_2_Z);
    
    \memory_memory_0_0_OLDA_RNIRSUT[6]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(6), C => 
        memory_memory_0_0_OLDA_Z(6), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(6));
    
    memoryrff_387_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya387_Z, B => WriteEnable, Y => 
        memorywre_387);
    
    memorya353_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(0), Y => memorya353_1_Z);
    
    memoryrff_494_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya494_Z, B => WriteEnable, Y => 
        memorywre_494);
    
    memoryrff_220_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya220_Z, B => WriteEnable, Y => 
        memorywre_220);
    
    memorya207 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya463_5_Z, B => memorya199_0_Z, C => 
        memorya482_2_Z, Y => memorya207_Z);
    
    \memory_memory_0_0_OLDA[3]\ : SLE
      port map(D => \InternalDataFromMem\(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(3));
    
    memoryrff_500 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_500, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_500);
    
    memoryrff_416 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_416, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_416);
    
    memorya54_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(4), Y => memorya54_2_Z);
    
    memory_memory_0_0_sr_RNO_379 : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory(3), B => memorya369_5_Z, 
        C => memorya441_6_Z, Y => memorya497);
    
    memory_memory_0_0_sr_RNO_45 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_133, B => memoryror_134, C => 
        memoryror_135, D => memoryror_132, Y => memoryror_417);
    
    memoryrff_96 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_96, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_96);
    
    memorya45_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya45_2_Z, B => memorya117_1_Z, Y => 
        memorya45_5_Z);
    
    memorya331_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya77_2_Z, B => memorya379_1_Z, Y => 
        memorya331_5_Z);
    
    memorya307 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya304_4_Z, 
        C => memorya379_4_Z, D => memorya499_5_Z, Y => 
        memorya307_Z);
    
    memory_memory_0_0_sr_RNO_218 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_435, B => memoryro_83, C => 
        memorya435, D => memorya83_Z, Y => memoryror_88);
    
    memoryrff_263_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya263_Z, B => WriteEnable, Y => 
        memorywre_263);
    
    memorya227_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya68_3_Z, B => InternalAddr2Memory(8), Y
         => memorya227_0_Z);
    
    memoryrff_108_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya108_Z, B => WriteEnable, Y => 
        memorywre_108);
    
    memoryrff_149 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_149, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_149);
    
    memoryrff_144_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya403_2_Z, B => WriteEnable, C => 
        memorya273_6_Z, D => memorya20_0_Z, Y => memorywre_144);
    
    memory_memory_0_0_sr_RNO_374 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya273_6_Z, B => memorya403_2_Z, C => 
        memorya20_0_Z, Y => memorya144);
    
    memoryrff_40 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_40, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_40);
    
    memorya276 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya84_3_Z, B => memorya273_4_Z, C => 
        memorya276_0_Z, D => memorya370_3_Z, Y => memorya276_Z);
    
    memoryrff_487_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya487_Z, B => WriteEnable, Y => 
        memorywre_487);
    
    memorya507 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya116_2_Z, B => InternalAddr2Memory(2), 
        C => memorya315_5_Z, D => memorya498_3_Z, Y => 
        memorya507_Z);
    
    memorya263 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya260_1_Z, B => memorya257_6_Z, C => 
        InternalAddr2Memory(7), D => memorya379_1_Z, Y => 
        memorya263_Z);
    
    memory_memory_0_0_sr_RNO_381 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya117_1_Z, B => memorya21_0_Z, C => 
        memorya20_6_Z, Y => memorya21);
    
    memorya233 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya233_0_Z, B => memorya121_1_Z, C => 
        memorya116_2_Z, D => memorya193_2_Z, Y => memorya233_Z);
    
    memory_memory_0_0_sr_RNO_239 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_87, B => memoryro_343, C => 
        memorya343_Z, D => memorya87_Z, Y => memoryror_78);
    
    memory_memory_0_0_sr_RNO_235 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_68, B => memoryro_468, C => 
        memorya468_Z, D => memorya68_Z, Y => memoryror_73);
    
    memoryrff_268 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_268, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_268);
    
    memorya280_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya125_2_Z, B => InternalAddr2Memory(7), 
        Y => memorya280_0_Z);
    
    memorya158 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya162_2_Z, B => memorya126_5_Z, C => 
        InternalAddr2Memory(8), D => memorya273_4_Z, Y => 
        memorya158_Z);
    
    memory_memory_0_0_sr_RNO_376 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya20_0_Z, B => memorya36_6_Z, C => 
        memorya36_1_Z, Y => memorya36);
    
    memoryrff_205 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_205, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_205);
    
    memoryrff_141_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya141_Z, B => WriteEnable, Y => 
        memorywre_141);
    
    memory_memory_0_0_sr_RNO_294 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_122, B => memoryro_506, C => 
        memorya506_Z, D => memorya122_Z, Y => memoryror_12);
    
    memoryrff_223_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya223_Z, B => WriteEnable, Y => 
        memorywre_223);
    
    memorya148 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya84_3_Z, B => memorya273_4_Z, C => 
        memorya52_0_Z, D => memorya162_2_Z, Y => memorya148_Z);
    
    \memory_memory_0_0_OLDA_RNI6IT31[10]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(10), C => 
        memory_memory_0_0_OLDA_Z(10), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(10));
    
    memoryrff_232 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_232, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_232);
    
    memory_memory_0_0_sr_RNO_302 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_379, B => memoryro_251, C => 
        memorya379_Z, D => memorya251, Y => memoryror_5);
    
    memoryrff_245_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya245_Z, B => WriteEnable, Y => 
        memorywre_245);
    
    memoryrff_145_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya145_Z, B => WriteEnable, Y => 
        memorywre_145);
    
    memorya65 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya57_3_Z, B => InternalAddr2Memory(8), C
         => memorya68_6_Z, D => memorya193_1_Z, Y => memorya65_Z);
    
    memorya47_0 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(4), Y => memorya47_0_Z);
    
    memorya364_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(2), Y => memorya364_1_Z);
    
    memory_memory_0_0_sr_RNO_195 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_354, B => memoryro_2, C => 
        memorya354_Z, D => memorya2_Z, Y => memoryror_128);
    
    \memory_memory_0_0_OLDA[25]\ : SLE
      port map(D => \InternalDataFromMem\(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(25));
    
    memorya112_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya54_2_Z, B => InternalAddr2Memory(8), Y
         => memorya63_0);
    
    memorya64 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya57_3_Z, B => InternalAddr2Memory(8), C
         => memorya68_6_Z, D => memorya84_2_Z, Y => memorya64_Z);
    
    \memory_memory_0_0_OLDA[0]\ : SLE
      port map(D => \InternalDataFromMem\(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(0));
    
    memoryrff_258_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya258_Z, B => WriteEnable, Y => 
        memorywre_258);
    
    memory_memory_0_0_sr_RNO_291 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_499, B => memoryro_51, C => 
        memorya499_Z, D => memorya51_Z, Y => memoryror_56);
    
    memoryrff_242_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya242_Z, B => WriteEnable, Y => 
        memorywre_242);
    
    memoryrff_238_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya238_Z, B => WriteEnable, Y => 
        memorywre_238);
    
    memory_memory_0_0_sr_RNO_317 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_41, B => memoryro_297, C => 
        memorya297_Z, D => memorya41_Z, Y => memoryror_45);
    
    memory_memory_0_0_sr_RNO_264 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_392, B => memoryro_8, C => 
        memorya392_Z, D => memorya8, Y => memoryror_127);
    
    memoryrff_79 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_79, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_79);
    
    memoryrff_388 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_388, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_388);
    
    \memory_memory_0_0_OLDA[1]\ : SLE
      port map(D => \InternalDataFromMem\(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(1));
    
    memoryrff_388_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya388_Z, B => WriteEnable, Y => 
        memorywre_388);
    
    memoryrff_350_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya350_Z, B => WriteEnable, Y => 
        memorywre_350);
    
    memorya286 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya273_4_Z, B => InternalAddr2Memory(7), 
        C => memorya126_5_Z, D => memorya370_3_Z, Y => 
        memorya286_Z);
    
    memory_memory_0_0_sr_RNO_359 : CFG3
      generic map(INIT => x"20")

      port map(A => memorya435_6_Z, B => InternalAddr2Memory(6), 
        C => memorya499_5_Z, Y => memorya435);
    
    memoryrff_415 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_415, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_415);
    
    memoryrff_330_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya330_Z, B => WriteEnable, Y => 
        memorywre_330);
    
    memoryrff_418_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya418_Z, B => WriteEnable, Y => 
        memorywre_418);
    
    memorya453 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya117_1_Z, B => InternalAddr2Memory(5), 
        C => memorya421_6_Z, D => memorya482_2_Z, Y => 
        memorya453_Z);
    
    memorya39 : CFG3
      generic map(INIT => x"20")

      port map(A => memorya36_6_Z, B => InternalAddr2Memory(8), C
         => memorya487_5_Z, Y => memorya39_Z);
    
    memorya8_0 : CFG3
      generic map(INIT => x"04")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(3), C => InternalAddr2Memory(8), Y
         => memorya8_0_Z);
    
    memorya152 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya56_0_Z, B => memorya162_2_Z, C => 
        memorya280_6_Z, Y => memorya152_Z);
    
    memory_memory_0_0_sr_RNO_320 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_293, B => memoryro_37, C => 
        memorya293, D => memorya37_Z, Y => memoryror_43);
    
    memory_memory_0_0_sr_RNO_290 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_52, B => memoryro_436, C => 
        memorya436_Z, D => memorya52_Z, Y => memoryror_57);
    
    memory_memory_0_0_sr_RNO_213 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_440, B => memoryro_40, C => 
        memorya440_Z, D => memorya40_Z, Y => memoryror_95);
    
    memorya443 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_4_Z, B => InternalAddr2Memory(6), 
        C => memorya315_5_Z, D => memorya434_2_Z, Y => 
        memorya443_Z);
    
    memorya40 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya52_4, B => memorya20_0_Z, C => 
        memorya41_3_Z, D => memorya45_2_Z, Y => memorya40_Z);
    
    memoryrff_406_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya406_Z, B => WriteEnable, Y => 
        memorywre_406);
    
    memorya142 : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory(8), B => memorya142_5_Z, 
        C => memorya270_6_Z, Y => memorya142_Z);
    
    memory_memory_0_0_sr_RNO_165 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_298, B => memoryro_154, C => 
        memorya298, D => memorya154_Z, Y => memoryror_156);
    
    memoryrff_293 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_293, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_293);
    
    memoryrff_194_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya194_Z, B => WriteEnable, Y => 
        memorywre_194);
    
    memorya84_2 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(0), Y => memorya84_2_Z);
    
    memorya301 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya289_4_Z, B => InternalAddr2Memory(7), 
        C => memorya45_5_Z, D => memorya369_3_Z, Y => 
        memorya301_Z);
    
    memorya142_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya395_2_Z, B => memorya102_1_Z, Y => 
        memorya142_5_Z);
    
    memory_memory_0_0_sr_RNO_365 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya503_5_Z, B => memorya111_0_Z, C => 
        memorya116_4_Z, Y => memorya119);
    
    memoryrff_211_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya211_Z, B => WriteEnable, Y => 
        memorywre_211);
    
    memory_memory_0_0_sr_RNO_261 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_382, B => memoryro_254, C => 
        memorya382_Z, D => memorya254_Z, Y => memoryror_119);
    
    \memory_memory_0_0_OLDA_RNIOPUT[3]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(3), C => 
        memory_memory_0_0_OLDA_Z(3), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(3));
    
    memoryrff_359_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya359_Z, B => WriteEnable, Y => 
        memorywre_359);
    
    memoryrff_302_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya302_Z, B => WriteEnable, Y => 
        memorywre_302);
    
    memoryrff_339_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya339_Z, B => WriteEnable, Y => 
        memorywre_339);
    
    memoryrff_449 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_449, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_449);
    
    memorya62 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya52_2_Z, C
         => memorya52_4, D => memorya126_5_Z, Y => memorya62_Z);
    
    memory_memory_0_0_sr_RNO_354 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya42_0_Z, B => memorya162_2_Z, C => 
        memorya264_6_Z, Y => memorya138);
    
    memory_memory_0_0_sr_RNO_24 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_227, B => memoryror_224, C => 
        memoryror_225, D => memoryror_226, Y => memoryror_440);
    
    memoryrff_10_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya362_1_Z, C => 
        memorya10_0_Z, D => memorya4_6_Z, Y => memorywre_10);
    
    memoryrff_191_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya191_Z, B => WriteEnable, Y => 
        memorywre_191);
    
    memory_memory_0_0_sr_RNO_260 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_125, B => memoryro_381, C => 
        memorya381_Z, D => memorya125_Z, Y => memoryror_118);
    
    memoryrff_313_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya313_Z, B => WriteEnable, Y => 
        memorywre_313);
    
    memorya257 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya257_0_Z, 
        C => memorya57_3_Z, D => memorya257_6_Z, Y => 
        memorya257_Z);
    
    memoryrff_488 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_488, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_488);
    
    memorya57 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya57_3_Z, C
         => memorya52_4, D => memorya121_5_Z, Y => memorya57_Z);
    
    memorya201 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya121_1_Z, 
        C => memorya393_6_Z, D => memorya482_2_Z, Y => 
        memorya201_Z);
    
    memory_memory_0_0_sr_RNO_356 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya9_0_Z, B => memorya264_6_Z, C => 
        memorya193_2_Z, Y => memorya137);
    
    memoryrff_93 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_93, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_93);
    
    memorya333_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya369_3_Z, B => memorya4_3_Z, Y => 
        memorya333_6_Z);
    
    memoryrff_295_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya295_Z, B => WriteEnable, Y => 
        memorywre_295);
    
    memorya436_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya434_2_Z, B => memorya116_1_Z, Y => 
        memorya436_5_Z);
    
    memorya423 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya68_3_Z, C
         => memorya487_5_Z, D => memorya498_3_Z, Y => 
        memorya423_Z);
    
    memoryrff_91_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya91_Z, B => WriteEnable, Y => 
        memorywre_91);
    
    memoryrff_31_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya31_Z, B => WriteEnable, Y => 
        memorywre_31);
    
    memoryrff_195_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya195_Z, B => WriteEnable, Y => 
        memorywre_195);
    
    memorya122 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya121_4_Z, 
        C => memorya84_2_Z, D => memorya378_5_Z, Y => 
        memorya122_Z);
    
    memoryrff_167 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_167, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_167);
    
    memorya357 : CFG3
      generic map(INIT => x"20")

      port map(A => memorya101_5_Z, B => InternalAddr2Memory(7), 
        C => memorya421_6_Z, Y => memorya357_Z);
    
    memoryrff_450_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya450_Z, B => WriteEnable, Y => 
        memorywre_450);
    
    memoryrff_292_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya292_Z, B => WriteEnable, Y => 
        memorywre_292);
    
    memoryrff_472_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya472_Z, B => WriteEnable, Y => 
        memorywre_472);
    
    memoryrff_430_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya430_Z, B => WriteEnable, Y => 
        memorywre_430);
    
    memorya87 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya68_4_Z, B => memorya503_5_Z, C => 
        memorya87_0, Y => memorya87_Z);
    
    \memory_memory_0_0_OLDA_RNIGTU31[29]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(29), C => 
        memory_memory_0_0_OLDA_Z(29), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(29));
    
    memorya347 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya25_3_Z, B => InternalAddr2Memory(7), C
         => memorya315_5_Z, D => memorya368_2_Z, Y => 
        memorya347_Z);
    
    memoryrff_152_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya152_Z, B => WriteEnable, Y => 
        memorywre_152);
    
    memoryrff_118 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_118, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_118);
    
    memoryrff_363 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_363, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_363);
    
    memoryrff_132_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya132_Z, B => WriteEnable, Y => 
        memorywre_132);
    
    memorya410 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya25_3_Z, B => InternalAddr2Memory(6), C
         => memorya154_5_Z, D => memorya370_3_Z, Y => 
        memorya410_Z);
    
    memorya492 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(4), B => memorya364_1_Z, 
        C => memorya116_2_Z, D => memorya504_6_Z, Y => 
        memorya492_Z);
    
    memoryrff_217 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_217, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_217);
    
    memoryrff_118_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya118_Z, B => WriteEnable, Y => 
        memorywre_118);
    
    memory_memory_0_0_sr_RNO_197 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_462, B => memoryro_62, C => 
        memorya462_Z, D => memorya62_Z, Y => memoryror_183);
    
    memoryrff_238 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_238, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_238);
    
    memorya227 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya211_3_Z, B => memorya379_1_Z, C => 
        memorya227_0_Z, D => memorya116_2_Z, Y => memorya227_Z);
    
    \memory_memory_0_0_OLDA[24]\ : SLE
      port map(D => \InternalDataFromMem\(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(24));
    
    memory_memory_0_0_sr_RNO_2 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_485, B => memoryror_484, C => 
        memoryror_486, D => memoryror_487, Y => memoryror_505);
    
    memorya7_0 : CFG2
      generic map(INIT => x"4")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(2), Y => memorya7_0_Z);
    
    memorya58 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya362_1_Z, B => memorya54_2_Z, C => 
        memorya52_4, D => memorya10_0_Z, Y => memorya58_Z);
    
    memoryrff_308 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_308, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_308);
    
    memorya264 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya68_2_Z, C
         => memorya264_1_Z, D => memorya264_6_Z, Y => 
        memorya264_Z);
    
    memorya234 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya233_0_Z, B => memorya362_1_Z, C => 
        memorya162_2_Z, D => memorya116_2_Z, Y => memorya234_Z);
    
    memory_memory_0_0_sr_RNO_328 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_363, B => memoryro_235, C => 
        memorya363_Z, D => memorya235_Z, Y => memoryror_21);
    
    memorya396 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya364_1_Z, 
        C => memorya204_6_Z, D => memorya498_3_Z, Y => 
        memorya396_Z);
    
    memorya327 : CFG3
      generic map(INIT => x"20")

      port map(A => memorya391_6_Z, B => InternalAddr2Memory(7), 
        C => memorya455_5_Z, Y => memorya327_Z);
    
    memory_memory_0_0_sr_RNO_209 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_307, B => memoryro_179, C => 
        memorya307_Z, D => memorya179_Z, Y => memoryror_184);
    
    memory_memory_0_0_sr_RNO_205 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_255, B => memoryro_447, C => 
        memorya447_Z, D => memorya255_Z, Y => memoryror_179);
    
    memoryrff_222 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_222, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_222);
    
    memorya79 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya79_0_Z, C
         => memorya463_5_Z, D => memorya68_4_Z, Y => memorya79_Z);
    
    memory_memory_0_0_sr_RNO_167 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_199, B => memoryro_407, C => 
        memorya407_Z, D => memorya199, Y => memoryror_158);
    
    \memory_memory_0_0_OLDA[20]\ : SLE
      port map(D => \InternalDataFromMem\(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(20));
    
    memory_memory_0_0_sr_RNO_133 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_368, B => memoryro_64, C => 
        memorya368, D => memorya64_Z, Y => memoryror_242);
    
    memoryrff_301_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya301_Z, B => WriteEnable, Y => 
        memorywre_301);
    
    memorya88 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya57_3_Z, B => memorya84_2_Z, C => 
        memorya56_0_Z, D => memorya68_4_Z, Y => memorya88_Z);
    
    memorya407 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya20_3_Z, C
         => memorya498_3_Z, D => memorya503_5_Z, Y => 
        memorya407_Z);
    
    memory_memory_0_0_sr_RNO_282 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_465, B => memoryro_113, C => 
        memorya465_Z, D => memorya113_Z, Y => memoryror_49);
    
    memoryrff_75 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_75, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_75);
    
    memorya506 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(2), B => memorya378_5_Z, 
        C => memorya370_3_Z, D => memorya482_2_Z, Y => 
        memorya506_Z);
    
    memorya295 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya289_4_Z, 
        C => memorya487_4_Z, D => memorya487_5_Z, Y => 
        memorya295_Z);
    
    memorya465 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya369_1_Z, B => InternalAddr2Memory(5), 
        C => memorya369_6_Z, D => memorya482_2_Z, Y => 
        memorya465_Z);
    
    memorya106 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya362_1_Z, B => memorya102_4_Z, C => 
        memorya116_2_Z, D => memorya10_0_Z, Y => memorya106_Z);
    
    memory_memory_0_0 : RAM1K18
      generic map(MEMORYFILE => "",
         RAMINDEX => "memory[31:0]%512-512%32-32%SPEED%0%0%TWO-PORT%ECC_EN-0"
        )

      port map(A_DOUT(17) => memory_memory_0_0_A_DOUT(17), 
        A_DOUT(16) => memory_memory_0_0_A_DOUT(16), A_DOUT(15)
         => memory_memory_0_0_A_DOUT(15), A_DOUT(14) => 
        memory_memory_0_0_A_DOUT(14), A_DOUT(13) => 
        memory_memory_0_0_NEWA(31), A_DOUT(12) => 
        memory_memory_0_0_NEWA(30), A_DOUT(11) => 
        memory_memory_0_0_NEWA(29), A_DOUT(10) => 
        memory_memory_0_0_NEWA(28), A_DOUT(9) => 
        memory_memory_0_0_NEWA(27), A_DOUT(8) => 
        memory_memory_0_0_NEWA(26), A_DOUT(7) => 
        memory_memory_0_0_NEWA(25), A_DOUT(6) => 
        memory_memory_0_0_NEWA(24), A_DOUT(5) => 
        memory_memory_0_0_NEWA(23), A_DOUT(4) => 
        memory_memory_0_0_NEWA(22), A_DOUT(3) => 
        memory_memory_0_0_NEWA(21), A_DOUT(2) => 
        memory_memory_0_0_NEWA(20), A_DOUT(1) => 
        memory_memory_0_0_NEWA(19), A_DOUT(0) => 
        memory_memory_0_0_NEWA(18), B_DOUT(17) => 
        memory_memory_0_0_NEWA(17), B_DOUT(16) => 
        memory_memory_0_0_NEWA(16), B_DOUT(15) => 
        memory_memory_0_0_NEWA(15), B_DOUT(14) => 
        memory_memory_0_0_NEWA(14), B_DOUT(13) => 
        memory_memory_0_0_NEWA(13), B_DOUT(12) => 
        memory_memory_0_0_NEWA(12), B_DOUT(11) => 
        memory_memory_0_0_NEWA(11), B_DOUT(10) => 
        memory_memory_0_0_NEWA(10), B_DOUT(9) => 
        memory_memory_0_0_NEWA(9), B_DOUT(8) => 
        memory_memory_0_0_NEWA(8), B_DOUT(7) => 
        memory_memory_0_0_NEWA(7), B_DOUT(6) => 
        memory_memory_0_0_NEWA(6), B_DOUT(5) => 
        memory_memory_0_0_NEWA(5), B_DOUT(4) => 
        memory_memory_0_0_NEWA(4), B_DOUT(3) => 
        memory_memory_0_0_NEWA(3), B_DOUT(2) => 
        memory_memory_0_0_NEWA(2), B_DOUT(1) => 
        memory_memory_0_0_NEWA(1), B_DOUT(0) => 
        memory_memory_0_0_NEWA(0), BUSY => NC0, A_CLK => 
        sb_sb_0_FIC_0_CLK, A_DOUT_CLK => \VCC\, A_ARST_N => \VCC\, 
        A_DOUT_EN => \VCC\, A_BLK(2) => \VCC\, A_BLK(1) => \VCC\, 
        A_BLK(0) => \VCC\, A_DOUT_ARST_N => \VCC\, A_DOUT_SRST_N
         => \VCC\, A_DIN(17) => \GND\, A_DIN(16) => \GND\, 
        A_DIN(15) => \GND\, A_DIN(14) => \GND\, A_DIN(13) => 
        InternalData2Memory(31), A_DIN(12) => 
        InternalData2Memory(30), A_DIN(11) => 
        InternalData2Memory(29), A_DIN(10) => 
        InternalData2Memory(28), A_DIN(9) => 
        InternalData2Memory(27), A_DIN(8) => 
        InternalData2Memory(26), A_DIN(7) => 
        InternalData2Memory(25), A_DIN(6) => 
        InternalData2Memory(24), A_DIN(5) => 
        InternalData2Memory(23), A_DIN(4) => 
        InternalData2Memory(22), A_DIN(3) => 
        InternalData2Memory(21), A_DIN(2) => 
        InternalData2Memory(20), A_DIN(1) => 
        InternalData2Memory(19), A_DIN(0) => 
        InternalData2Memory(18), A_ADDR(13) => 
        InternalAddr2Memory(8), A_ADDR(12) => 
        InternalAddr2Memory(7), A_ADDR(11) => 
        InternalAddr2Memory(6), A_ADDR(10) => 
        InternalAddr2Memory(5), A_ADDR(9) => 
        InternalAddr2Memory(4), A_ADDR(8) => 
        InternalAddr2Memory(3), A_ADDR(7) => 
        InternalAddr2Memory(2), A_ADDR(6) => 
        InternalAddr2Memory(1), A_ADDR(5) => 
        InternalAddr2Memory(0), A_ADDR(4) => \GND\, A_ADDR(3) => 
        \GND\, A_ADDR(2) => \GND\, A_ADDR(1) => \GND\, A_ADDR(0)
         => \GND\, A_WEN(1) => \VCC\, A_WEN(0) => \VCC\, B_CLK
         => sb_sb_0_FIC_0_CLK, B_DOUT_CLK => \VCC\, B_ARST_N => 
        \VCC\, B_DOUT_EN => \VCC\, B_BLK(2) => WriteEnable, 
        B_BLK(1) => WriteEnable, B_BLK(0) => WriteEnable, 
        B_DOUT_ARST_N => \VCC\, B_DOUT_SRST_N => \VCC\, B_DIN(17)
         => InternalData2Memory(17), B_DIN(16) => 
        InternalData2Memory(16), B_DIN(15) => 
        InternalData2Memory(15), B_DIN(14) => 
        InternalData2Memory(14), B_DIN(13) => 
        InternalData2Memory(13), B_DIN(12) => 
        InternalData2Memory(12), B_DIN(11) => 
        InternalData2Memory(11), B_DIN(10) => 
        InternalData2Memory(10), B_DIN(9) => 
        InternalData2Memory(9), B_DIN(8) => 
        InternalData2Memory(8), B_DIN(7) => 
        InternalData2Memory(7), B_DIN(6) => 
        InternalData2Memory(6), B_DIN(5) => 
        InternalData2Memory(5), B_DIN(4) => 
        InternalData2Memory(4), B_DIN(3) => 
        InternalData2Memory(3), B_DIN(2) => 
        InternalData2Memory(2), B_DIN(1) => 
        InternalData2Memory(1), B_DIN(0) => 
        InternalData2Memory(0), B_ADDR(13) => 
        InternalAddr2Memory(8), B_ADDR(12) => 
        InternalAddr2Memory(7), B_ADDR(11) => 
        InternalAddr2Memory(6), B_ADDR(10) => 
        InternalAddr2Memory(5), B_ADDR(9) => 
        InternalAddr2Memory(4), B_ADDR(8) => 
        InternalAddr2Memory(3), B_ADDR(7) => 
        InternalAddr2Memory(2), B_ADDR(6) => 
        InternalAddr2Memory(1), B_ADDR(5) => 
        InternalAddr2Memory(0), B_ADDR(4) => \GND\, B_ADDR(3) => 
        \GND\, B_ADDR(2) => \GND\, B_ADDR(1) => \GND\, B_ADDR(0)
         => \GND\, B_WEN(1) => \VCC\, B_WEN(0) => \VCC\, A_EN => 
        \VCC\, A_DOUT_LAT => \VCC\, A_WIDTH(2) => \VCC\, 
        A_WIDTH(1) => \VCC\, A_WIDTH(0) => \GND\, A_WMODE => 
        \GND\, B_EN => \VCC\, B_DOUT_LAT => \VCC\, B_WIDTH(2) => 
        \VCC\, B_WIDTH(1) => \VCC\, B_WIDTH(0) => \GND\, B_WMODE
         => \GND\, SII_LOCK => \GND\);
    
    memorya432_0 : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory(6), B => memorya54_2_Z, C
         => memorya498_3_Z, Y => memorya432_0_Z);
    
    memoryrff_77 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_77, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_77);
    
    memoryrff_246_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya246_Z, B => WriteEnable, Y => 
        memorywre_246);
    
    memorya45 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya45_2_Z, B => memorya45_6_Z, C => 
        InternalAddr2Memory(8), D => memorya117_1_Z, Y => 
        memorya45_Z);
    
    memoryrff_253 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_253, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_253);
    
    memorya373_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya54_2_Z, B => memorya117_1_Z, Y => 
        memorya373_5_Z);
    
    memoryrff_408 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_408, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_408);
    
    memorya351 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya415_4_Z, 
        C => memorya86_2_Z, D => memorya463_5_Z, Y => 
        memorya351_Z);
    
    memorya100 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya36_1_Z, C
         => memorya84_2_Z, D => memorya100_6_Z, Y => memorya100_Z);
    
    \memory_memory_0_0_OLDA_RNI9NV31[31]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(31), C => 
        memory_memory_0_0_OLDA_Z(31), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(31));
    
    memoryrff_416_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya416_Z, B => WriteEnable, Y => 
        memorywre_416);
    
    memoryrff_273 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_273, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_273);
    
    memorya341 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya20_3_Z, B => InternalAddr2Memory(7), C
         => memorya213_5_Z, D => memorya369_3_Z, Y => 
        memorya341_Z);
    
    memorya193 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya193_1_Z, 
        C => memorya193_2_Z, D => memorya320_6_Z, Y => 
        memorya193_Z);
    
    memoryrff_453_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya453_Z, B => WriteEnable, Y => 
        memorywre_453);
    
    memoryrff_433_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya433_Z, B => WriteEnable, Y => 
        memorywre_433);
    
    memoryrff_312_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya312_Z, B => WriteEnable, Y => 
        memorywre_312);
    
    memorya296_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya289_4_Z, B => memorya57_3_Z, Y => 
        memorya296_6_Z);
    
    memory_memory_0_0_sr_RNO_41 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_149, B => memoryror_151, C => 
        memoryror_148, D => memoryror_150, Y => memoryror_421);
    
    memoryrff_137 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_137, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_137);
    
    memoryrff_92 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_92, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_92);
    
    memoryrff_376_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya376_Z, B => WriteEnable, Y => 
        memorywre_376);
    
    memoryrff_361 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_361, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_361);
    
    memorya318_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(0), Y => memorya318_4_Z);
    
    memorya42 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya41_3_Z, B => memorya52_2_Z, C => 
        memorya42_0_Z, D => memorya52_4, Y => memorya42_Z);
    
    memorya321 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya193_1_Z, B => InternalAddr2Memory(7), 
        C => memorya320_6_Z, D => memorya369_3_Z, Y => 
        memorya321_Z);
    
    memoryrff_333 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_333, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_333);
    
    memoryrff_165 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_165, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_165);
    
    memoryrff_314 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_314, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_314);
    
    memorya369_3 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(1), Y => memorya369_3_Z);
    
    memory_memory_0_0_sr_RNO_191 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_169, B => memoryro_409, C => 
        memorya409_Z, D => memorya169_Z, Y => memoryror_141);
    
    memory_memory_0_0_sr_RNO_124 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_463, B => memoryro_143, C => 
        memorya463_Z, D => memorya143_Z, Y => memoryror_195);
    
    memory_memory_0_0_sr_RNO_237 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_56, B => memoryro_424, C => 
        memorya424_Z, D => memorya56_Z, Y => memoryror_79);
    
    memoryrff_296_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya296_Z, B => WriteEnable, Y => 
        memorywre_296);
    
    memorya455_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya68_1_Z, B => memorya379_1_Z, Y => 
        memorya455_5_Z);
    
    memorya177 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya369_1_Z, B => InternalAddr2Memory(8), 
        C => memorya304_6_Z, D => memorya434_2_Z, Y => 
        memorya177_Z);
    
    memoryrff_228 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_228, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_228);
    
    memoryrff_289 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_289, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_289);
    
    memorya221 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya29_3_Z, C
         => memorya381_5_Z, D => memorya482_2_Z, Y => 
        memorya221_Z);
    
    memoryrff_180_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya180_Z, B => WriteEnable, Y => 
        memorywre_180);
    
    memorya86_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(4), Y => memorya86_2_Z);
    
    memory_memory_0_0_sr_RNO_161 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_445, B => memoryro_221, C => 
        memorya445_Z, D => memorya221_Z, Y => memoryror_166);
    
    memorya11_0 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(2), Y => memorya11_0_Z);
    
    memorya116_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(5), Y => memorya116_2_Z);
    
    memoryrff_186 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_186, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_186);
    
    memory_memory_0_0_sr_RNO_319 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_90, B => memoryro_474, C => 
        memorya474_Z, D => memorya90_Z, Y => memoryror_44);
    
    memoryrff_146_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya146_Z, B => WriteEnable, Y => 
        memorywre_146);
    
    memorya457 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya121_1_Z, B => InternalAddr2Memory(5), 
        C => memorya361_6_Z, D => memorya482_2_Z, Y => 
        memorya457_Z);
    
    \memory_memory_0_0_OLDA_RNIDQU31[26]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(26), C => 
        memory_memory_0_0_OLDA_Z(26), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(26));
    
    memoryrff_292 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_292, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_292);
    
    memorya447 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya364_1_Z, B => memorya432_0_Z, C => 
        InternalAddr2Memory(1), D => InternalAddr2Memory(0), Y
         => memorya447_Z);
    
    memory_memory_0_0_sr_RNO_284 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_203, B => memoryro_331, C => 
        memorya331_Z, D => memorya203, Y => memoryror_53);
    
    memoryrff_489_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya489_Z, B => WriteEnable, Y => 
        memorywre_489);
    
    memoryrff_311_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya311_Z, B => WriteEnable, Y => 
        memorywre_311);
    
    memorya296 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya45_2_Z, B => InternalAddr2Memory(7), C
         => memorya296_6_Z, D => memorya370_3_Z, Y => 
        memorya296_Z);
    
    memory_memory_0_0_sr_RNO_103 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_352, B => memoryro_80, C => 
        memorya352_Z, D => memorya80, Y => memoryror_226);
    
    memorya156 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_2_Z, B => InternalAddr2Memory(8), C
         => memorya156_5_Z, D => memorya273_4_Z, Y => 
        memorya156_Z);
    
    memoryrff_463 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_463, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_463);
    
    memoryrff_460 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_460, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_460);
    
    memorya187 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya312_4_Z, B => InternalAddr2Memory(8), 
        C => memorya315_5_Z, D => memorya434_2_Z, Y => 
        memorya187_Z);
    
    memorya372 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya116_1_Z, 
        C => memorya116_2_Z, D => memorya372_6_Z, Y => 
        memorya372_Z);
    
    memorya146 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya162_2_Z, B => memorya273_6_Z, C => 
        InternalAddr2Memory(8), D => memorya370_1_Z, Y => 
        memorya146_Z);
    
    memoryrff_204_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya204_Z, B => WriteEnable, Y => 
        memorywre_204);
    
    memorya179 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya304_4_Z, 
        C => memorya211_3_Z, D => memorya499_5_Z, Y => 
        memorya179_Z);
    
    memory_memory_0_0_sr_RNO_176 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_145, B => memoryro_273, C => 
        memorya273_Z, D => memorya145_Z, Y => memoryror_145);
    
    memory_memory_0_0_sr_RNO_314 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_449, B => memoryro_97, C => 
        memorya449_Z, D => memorya97_Z, Y => memoryror_33);
    
    memory_memory_0_0_sr_RNO_185 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_413, B => memoryro_253, C => 
        memorya413_Z, D => memorya253_Z, Y => memoryror_134);
    
    memoryrff_83_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya83_Z, B => WriteEnable, Y => 
        memorywre_83);
    
    memoryrff_66 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_66, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_66);
    
    memoryrff_458_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya458_Z, B => WriteEnable, Y => 
        memorywre_458);
    
    memoryrff_438_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya438_Z, B => WriteEnable, Y => 
        memorywre_438);
    
    memorya150 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_1_Z, B => InternalAddr2Memory(8), 
        C => memorya278_6_Z, D => memorya403_2_Z, Y => 
        memorya150_Z);
    
    memorya118 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya84_2_Z, C
         => memorya116_4_Z, D => memorya118_5_Z, Y => 
        memorya118_Z);
    
    memory_memory_0_0_sr_RNO_281 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_496, B => memoryro_128, C => 
        memorya496_Z, D => memorya128, Y => memoryror_50);
    
    memoryrff_74 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_74, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_74);
    
    memorya140 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya12_0_Z, B => memorya162_2_Z, C => 
        memorya268_6_Z, Y => memorya140_Z);
    
    memoryrff_164 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_164, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_164);
    
    memorya479 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya364_1_Z, B => memorya464_0_Z, C => 
        InternalAddr2Memory(1), D => InternalAddr2Memory(0), Y
         => memorya479_Z);
    
    memorya373 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya84_3_Z, C
         => memorya368_2_Z, D => memorya373_5_Z, Y => 
        memorya373_Z);
    
    memory_memory_0_0_sr_RNO_316 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_88, B => memoryro_488, C => 
        memorya488_Z, D => memorya88_Z, Y => memoryror_47);
    
    memoryrff_251_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya211_3_Z, C => 
        memorya315_5_Z, D => memorya111_0_Z, Y => memorywre_251);
    
    memorya427 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya41_3_Z, B => InternalAddr2Memory(6), C
         => memorya299_5_Z, D => memorya498_3_Z, Y => 
        memorya427_Z);
    
    memoryrff_231_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya231_Z, B => WriteEnable, Y => 
        memorywre_231);
    
    memorya4_0 : CFG2
      generic map(INIT => x"4")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(2), Y => memorya4_0_Z);
    
    memorya204_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya4_3_Z, B => memorya68_2_Z, Y => 
        memorya204_6_Z);
    
    memory_memory_0_0_sr_RNO_280 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_63, B => memoryro_319, C => 
        memorya319_Z, D => memorya63_Z, Y => memoryror_51);
    
    \memory_memory_0_0_OLDA_RNI8MV31[30]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(30), C => 
        memory_memory_0_0_OLDA_Z(30), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(30));
    
    memoryrff_189_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya189_Z, B => WriteEnable, Y => 
        memorywre_189);
    
    memorya61 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya37_2_Z, C
         => memorya52_4, D => memorya381_5_Z, Y => memorya61_Z);
    
    memorya161 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya193_2_Z, B => memorya289_6_Z, C => 
        InternalAddr2Memory(8), D => memorya353_1_Z, Y => 
        memorya161_Z);
    
    memoryrff_331 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_331, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_331);
    
    memoryrff_110 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_110, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_110);
    
    memoryrff_462_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya462_Z, B => WriteEnable, Y => 
        memorywre_462);
    
    memoryrff_243 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_243, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_243);
    
    memorya131 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya211_3_Z, B => memorya257_6_Z, C => 
        InternalAddr2Memory(8), D => memorya379_1_Z, Y => 
        memorya131_Z);
    
    memorya126 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya126_0_Z, 
        C => memorya116_2_Z, D => memorya126_5_Z, Y => 
        memorya126_Z);
    
    memoryrff_58 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_58, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_58);
    
    memoryrff_353_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya353_Z, B => WriteEnable, Y => 
        memorywre_353);
    
    memoryrff_127 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_127, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_127);
    
    memoryrff_387 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_387, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_387);
    
    memoryrff_36 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_36, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_36);
    
    memoryrff_333_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya333_Z, B => WriteEnable, Y => 
        memorywre_333);
    
    memorya498_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya498_3_Z, B => memorya354_3_Z, Y => 
        memorya498_6_Z);
    
    memoryrff_196_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya196_Z, B => WriteEnable, Y => 
        memorywre_196);
    
    memoryrff_135 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_135, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_135);
    
    memorya382 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya116_2_Z, B => InternalAddr2Memory(7), 
        C => memorya126_5_Z, D => memorya370_3_Z, Y => 
        memorya382_Z);
    
    memoryrff_99 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_99, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_99);
    
    memorya413 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya29_3_Z, B => InternalAddr2Memory(6), C
         => memorya381_5_Z, D => memorya498_3_Z, Y => 
        memorya413_Z);
    
    memorya189 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya316_4_Z, B => InternalAddr2Memory(8), 
        C => memorya381_5_Z, D => memorya434_2_Z, Y => 
        memorya189_Z);
    
    memorya112 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya84_2_Z, B => memorya57_3_Z, C => 
        memorya63_0, D => memorya116_4_Z, Y => memorya112_Z);
    
    memory_memory_0_0_sr_RNO_362 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya111_0_Z, B => memorya102_4_Z, C => 
        memorya463_5_Z, Y => memorya111);
    
    memory_memory_0_0_sr_RNO_178 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_272, B => memoryro_32, C => 
        memorya272_Z, D => memorya32_Z, Y => memoryror_146);
    
    memoryrff_209 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_209, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_209);
    
    memorya120 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya125_2_Z, B => memorya121_4_Z, C => 
        memorya116_2_Z, D => memorya20_0_Z, Y => memorya120_Z);
    
    memoryrff_323 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_323, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_323);
    
    memoryrff_441_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya441_Z, B => WriteEnable, Y => 
        memorywre_441);
    
    memorya360 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya45_2_Z, C
         => memorya360_6_Z, D => memorya368_2_Z, Y => 
        memorya360_Z);
    
    memorya330 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya202_6_Z, B => memorya368_2_Z, C => 
        memorya266_0_Z, Y => memorya330_Z);
    
    memorya489 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(4), B => memorya121_1_Z, 
        C => memorya116_2_Z, D => memorya441_6_Z, Y => 
        memorya489_Z);
    
    memorya383 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya364_1_Z, B => memorya368_0_Z, C => 
        InternalAddr2Memory(1), D => InternalAddr2Memory(0), Y
         => memorya383_Z);
    
    memoryrff_79_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya79_Z, B => WriteEnable, Y => 
        memorywre_79);
    
    memoryrff_422_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya422_Z, B => WriteEnable, Y => 
        memorywre_422);
    
    memorya10_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya354_3_Z, B => InternalAddr2Memory(8), 
        Y => memorya10_0_Z);
    
    memorya104 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya45_2_Z, C
         => memorya84_2_Z, D => memorya105_6_Z, Y => memorya104_Z);
    
    memoryrff_278_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya278_Z, B => WriteEnable, Y => 
        memorywre_278);
    
    memoryrff_106 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_106, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_106);
    
    memorya59 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya35_0_Z, B => memorya52_4, C => 
        memorya315_5_Z, Y => memorya59_Z);
    
    memory_memory_0_0_sr_RNO_156 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_423, B => memoryro_247, C => 
        memorya423_Z, D => memorya247, Y => memoryror_174);
    
    memoryrff_404_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya404_Z, B => WriteEnable, Y => 
        memorywre_404);
    
    memory_memory_0_0_sr_RNO_207 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_305, B => memoryro_177, C => 
        memorya305_Z, D => memorya177_Z, Y => memoryror_177);
    
    \memory_memory_0_0_OLDA_RNI9LT31[13]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(13), C => 
        memory_memory_0_0_OLDA_Z(13), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(13));
    
    memoryrff_158_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya158_Z, B => WriteEnable, Y => 
        memorywre_158);
    
    memorya217 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya25_3_Z, C
         => memorya193_2_Z, D => memorya345_5_Z, Y => 
        memorya217_Z);
    
    memoryrff_370_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya370_Z, B => WriteEnable, Y => 
        memorywre_370);
    
    memoryrff_298 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_298, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_298);
    
    memoryrff_138_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya162_2_Z, B => memorya264_6_Z, C => 
        WriteEnable, D => memorya42_0_Z, Y => memorywre_138);
    
    memory_memory_0_0_sr_RNO_22 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_216, B => memoryror_219, C => 
        memoryror_217, D => memoryror_218, Y => memoryror_438);
    
    memoryrff_266 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_266, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_266);
    
    memory_memory_0_0_sr_RNO_53 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_91, B => memoryror_89, C => 
        memoryror_88, D => memoryror_90, Y => memoryror_406);
    
    memory_memory_0_0_sr_RNO_74 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_6, B => memoryror_7, C => 
        memoryror_5, D => memoryror_4, Y => memoryror_385);
    
    memory_memory_0_0_sr_RNO_187 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_332, B => memoryro_140, C => 
        memorya332_Z, D => memorya140_Z, Y => memoryror_132);
    
    memorya89 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya57_3_Z, C
         => memorya68_4_Z, D => memorya345_5_Z, Y => memorya89_Z);
    
    memorya317 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya316_4_Z, 
        C => memorya305_2_Z, D => memorya381_5_Z, Y => 
        memorya317_Z);
    
    memoryrff_379_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya379_Z, B => WriteEnable, Y => 
        memorywre_379);
    
    memoryrff_252 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_252, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_252);
    
    memorya468 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya116_1_Z, B => InternalAddr2Memory(5), 
        C => memorya372_6_Z, D => memorya482_2_Z, Y => 
        memorya468_Z);
    
    memorya364 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya364_1_Z, 
        C => memorya116_2_Z, D => memorya364_6_Z, Y => 
        memorya364_Z);
    
    memoryrff_72_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya72_Z, B => WriteEnable, Y => 
        memorywre_72);
    
    memoryrff_433 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_433, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_433);
    
    memoryrff_430 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_430, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_430);
    
    memoryrff_272 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_272, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_272);
    
    memorya438 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_3_Z, B => InternalAddr2Memory(6), 
        C => memorya118_5_Z, D => memorya498_3_Z, Y => 
        memorya438_Z);
    
    memorya334 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya4_3_Z, B => InternalAddr2Memory(7), C
         => memorya78_5_Z, D => memorya370_3_Z, Y => memorya334_Z);
    
    memorya126_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya102_1_Z, B => memorya125_2_Z, Y => 
        memorya126_5_Z);
    
    memoryrff_183 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_183, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_183);
    
    memorya19_0 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(2), Y => memorya19_0_Z);
    
    memory_memory_0_0_sr_RNO_83 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_27, B => memoryror_24, C => 
        memoryror_26, D => memoryror_25, Y => memoryror_390);
    
    memorya404 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya116_1_Z, 
        C => memorya340_6_Z, D => memorya498_3_Z, Y => 
        memorya404_Z);
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    memory_memory_0_0_sr_RNO_333 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_25, B => memoryro_281, C => 
        memorya281_Z, D => memorya25_Z, Y => memoryror_29);
    
    memoryrff_63 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_63, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_63);
    
    memoryrff_491_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya491_Z, B => WriteEnable, Y => 
        memorywre_491);
    
    memory_memory_0_0_sr_RNO_158 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_216, B => memoryro_296, C => 
        memorya296_Z, D => memorya216_Z, Y => memoryror_175);
    
    memory_memory_0_0_sr_RNO_17 : CFG4
      generic map(INIT => x"0001")

      port map(A => memoryror_387, B => memoryror_386, C => 
        memoryror_385, D => memoryror_384, Y => memoryror_504_1);
    
    memoryrff_134 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_134, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_134);
    
    memorya165 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya117_1_Z, B => InternalAddr2Memory(8), 
        C => memorya292_6_Z, D => memorya434_2_Z, Y => 
        memorya165_Z);
    
    \memory_memory_0_0_OLDA[8]\ : SLE
      port map(D => \InternalDataFromMem\(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(8));
    
    memoryrff_6_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya6_Z, B => WriteEnable, Y => 
        memorywre_6);
    
    memoryrff_214_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya214_Z, B => WriteEnable, Y => 
        memorywre_214);
    
    memoryrff_50 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_50, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_50);
    
    memorya135 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_1_Z, B => InternalAddr2Memory(8), 
        C => memorya257_6_Z, D => memorya391_2_Z, Y => 
        memorya135_Z);
    
    memoryrff_347_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya347_Z, B => WriteEnable, Y => 
        memorywre_347);
    
    memoryrff_307 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_307, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_307);
    
    memorya395_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya395_2_Z, B => memorya379_1_Z, Y => 
        memorya395_5_Z);
    
    memorya213_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya86_2_Z, B => memorya117_1_Z, Y => 
        memorya213_5_Z);
    
    memoryrff_84_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya84_Z, B => WriteEnable, Y => 
        memorywre_84);
    
    memoryrff_470_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya470_Z, B => WriteEnable, Y => 
        memorywre_470);
    
    memoryrff_366_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya366_Z, B => WriteEnable, Y => 
        memorywre_366);
    
    memory_memory_0_0_sr_RNO_299 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_3, B => memoryro_451, C => 
        memorya451_Z, D => memorya3, Y => memoryror_8);
    
    memory_memory_0_0_sr_RNO_295 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_456, B => memoryro_120, C => 
        memorya456_Z, D => memorya120_Z, Y => memoryror_15);
    
    memoryrff_456_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya456_Z, B => WriteEnable, Y => 
        memorywre_456);
    
    memoryrff_436_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya436_Z, B => WriteEnable, Y => 
        memorywre_436);
    
    memoryrff_172_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya172_Z, B => WriteEnable, Y => 
        memorywre_172);
    
    memorya110_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya45_2_Z, B => memorya102_1_Z, Y => 
        memorya110_5_Z);
    
    memory_memory_0_0_sr_RNO_7 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_444, B => memoryror_447, C => 
        memoryror_445, D => memoryror_446, Y => memoryror_495);
    
    memoryrff_33 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_33, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_33);
    
    memoryrff_352_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya352_Z, B => WriteEnable, Y => 
        memorywre_352);
    
    memoryrff_332_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya332_Z, B => WriteEnable, Y => 
        memorywre_332);
    
    memoryrff_321 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_321, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_321);
    
    memory_memory_0_0_sr_RNO_246 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_58, B => memoryro_442, C => 
        memorya442_Z, D => memorya58_Z, Y => memoryror_108);
    
    memoryrff_161 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_161, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_161);
    
    \memory_memory_0_0_OLDA_RNIMNUT[1]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(1), C => 
        memory_memory_0_0_OLDA_Z(1), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(1));
    
    memoryrff_95 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_95, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_95);
    
    memoryrff_197 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_197, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_197);
    
    memoryrff_125 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_125, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_125);
    
    memory_memory_0_0_sr_RNO_269 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_242, B => memoryro_402, C => 
        memorya402_Z, D => memorya242_Z, Y => memoryror_112);
    
    memory_memory_0_0_sr_RNO_265 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_377, B => memoryro_121, C => 
        memorya377_Z, D => memorya121_Z, Y => memoryror_125);
    
    memoryrff_97 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_97, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_97);
    
    memoryrff_326_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya326_Z, B => WriteEnable, Y => 
        memorywre_326);
    
    memorya41 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya52_4, B => memorya9_0_Z, C => 
        memorya37_2_Z, D => memorya41_3_Z, Y => memorya41_Z);
    
    memoryrff_90_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya90_Z, B => WriteEnable, Y => 
        memorywre_90);
    
    memoryrff_30_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya30_Z, B => WriteEnable, Y => 
        memorywre_30);
    
    memorya311 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya304_4_Z, 
        C => memorya305_2_Z, D => memorya503_5_Z, Y => 
        memorya311_Z);
    
    memoryrff_43_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya43_Z, B => WriteEnable, Y => 
        memorywre_43);
    
    memoryrff_104_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya104_Z, B => WriteEnable, Y => 
        memorywre_104);
    
    memoryrff_393 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_393, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_393);
    
    memoryrff_466 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_466, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_466);
    
    memoryrff_1 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_1, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_1);
    
    memoryrff_447_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya447_Z, B => WriteEnable, Y => 
        memorywre_447);
    
    memorya154 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya273_4_Z, B => memorya154_5_Z, C => 
        InternalAddr2Memory(8), D => memorya354_3_Z, Y => 
        memorya154_Z);
    
    memoryrff_236 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_236, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_236);
    
    memorya375 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya487_4_Z, 
        C => memorya116_2_Z, D => memorya503_5_Z, Y => 
        memorya375_Z);
    
    memorya309 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya304_4_Z, 
        C => memorya369_3_Z, D => memorya373_5_Z, Y => 
        memorya309_Z);
    
    memoryrff_397_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya397_Z, B => WriteEnable, Y => 
        memorywre_397);
    
    memoryrff_101_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya101_Z, B => WriteEnable, Y => 
        memorywre_101);
    
    memoryrff_258 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_258, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_258);
    
    memorya435_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya498_3_Z, B => memorya368_4_Z, Y => 
        memorya435_6_Z);
    
    memorya239 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya116_2_Z, B => memorya463_5_Z, C => 
        memorya143_0_Z, Y => memorya239_Z);
    
    memory_memory_0_0_sr_RNO_181 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_181, B => memoryro_405, C => 
        memorya405_Z, D => memorya181_Z, Y => memoryror_139);
    
    memory_memory_0_0_sr_RNO_15 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_413, B => memoryror_415, C => 
        memoryror_412, D => memoryror_414, Y => memoryror_487);
    
    memorya211 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya211_3_Z, B => memorya211_0_Z, C => 
        memorya379_1_Z, D => memorya86_2_Z, Y => memorya211_Z);
    
    memoryrff_414_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya414_Z, B => WriteEnable, Y => 
        memorywre_414);
    
    memorya362_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya370_3_Z, B => memorya41_3_Z, Y => 
        memorya362_6_Z);
    
    memoryrff_278 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_278, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_278);
    
    memoryrff_205_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya205_Z, B => WriteEnable, Y => 
        memorywre_205);
    
    memoryrff_103 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_103, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_103);
    
    memoryrff_7_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya7_Z, B => WriteEnable, Y => 
        memorywre_7);
    
    memoryrff_105_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya105_Z, B => WriteEnable, Y => 
        memorywre_105);
    
    memory_memory_0_0_sr_RNO_50 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_176, B => memoryror_179, C => 
        memoryror_178, D => memoryror_177, Y => memoryror_428);
    
    memory_memory_0_0_sr_RNO_179 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_18, B => memoryro_370, C => 
        memorya370_Z, D => memorya18, Y => memoryror_144);
    
    memoryrff_189 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_189, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_189);
    
    memorya463_5 : CFG3
      generic map(INIT => x"80")

      port map(A => InternalAddr2Memory(0), B => memorya364_1_Z, 
        C => InternalAddr2Memory(1), Y => memorya463_5_Z);
    
    memory_memory_0_0_sr_RNO_170 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_348, B => memoryro_156, C => 
        memorya348_Z, D => memorya156_Z, Y => memoryror_148);
    
    memorya466 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya370_1_Z, B => InternalAddr2Memory(5), 
        C => memorya370_6_Z, D => memorya482_2_Z, Y => 
        memorya466_Z);
    
    memorya403_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(4), Y => memorya403_2_Z);
    
    memoryrff_348_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya348_Z, B => WriteEnable, Y => 
        memorywre_348);
    
    memoryrff_202_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya202_Z, B => WriteEnable, Y => 
        memorywre_202);
    
    memorya436 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya116_1_Z, B => InternalAddr2Memory(6), 
        C => memorya372_6_Z, D => memorya434_2_Z, Y => 
        memorya436_Z);
    
    memoryrff_411 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_411, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_411);
    
    memoryrff_473_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya473_Z, B => WriteEnable, Y => 
        memorywre_473);
    
    memoryrff_423 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_423, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_423);
    
    memoryrff_420 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_420, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_420);
    
    memoryrff_8 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_8, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_8);
    
    memorya197 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya117_1_Z, 
        C => memorya197_6_Z, D => memorya482_2_Z, Y => 
        memorya197_Z);
    
    memoryrff_211 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_211, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_211);
    
    memory_memory_0_0_sr_RNO_330 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_124, B => memoryro_396, C => 
        memorya396_Z, D => memorya124, Y => memoryror_20);
    
    memoryrff_485_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya485_Z, B => WriteEnable, Y => 
        memorywre_485);
    
    memoryrff_351_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya351_Z, B => WriteEnable, Y => 
        memorywre_351);
    
    memoryrff_2_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya2_Z, B => WriteEnable, Y => 
        memorywre_2);
    
    memorya454 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_1_Z, B => InternalAddr2Memory(5), 
        C => memorya358_6_Z, D => memorya482_2_Z, Y => 
        memorya454_Z);
    
    memorya17 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya57_3_Z, B => memorya20_6_Z, C => 
        InternalAddr2Memory(8), D => memorya369_1_Z, Y => 
        memorya17_Z);
    
    \memory_memory_0_0_OLDA_RNI7JT31[11]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(11), C => 
        memory_memory_0_0_OLDA_Z(11), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(11));
    
    memoryrff_331_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya331_Z, B => WriteEnable, Y => 
        memorywre_331);
    
    memoryrff_62 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_62, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_62);
    
    memoryrff_19_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya19_Z, B => WriteEnable, Y => 
        memorywre_19);
    
    memorya385 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya369_3_Z, B => memorya320_6_Z, C => 
        InternalAddr2Memory(6), D => memorya385_1_Z, Y => 
        memorya385_Z);
    
    memorya444 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_2_Z, B => InternalAddr2Memory(6), C
         => memorya380_5_Z, D => memorya498_3_Z, Y => 
        memorya444_Z);
    
    memory_memory_0_0_sr_RNO_64 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_118, B => memoryror_119, C => 
        memoryror_116, D => memoryror_117, Y => memoryror_413);
    
    \memory_memory_0_0_OLDA[26]\ : SLE
      port map(D => \InternalDataFromMem\(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(26));
    
    memoryrff_242 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_242, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_242);
    
    memorya101_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya116_2_Z, B => memorya117_1_Z, Y => 
        memorya101_5_Z);
    
    memory_memory_0_0_sr_RNO_80 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_19, B => memoryror_18, C => 
        memoryror_17, D => memoryror_16, Y => memoryror_388);
    
    memoryrff_497_RNO : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya369_5_Z, B => memorya441_6_Z, C => 
        InternalAddr2Memory(3), D => WriteEnable, Y => 
        memorywre_497);
    
    memorya4_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(4), Y => memorya4_3_Z);
    
    memory_memory_0_0_sr_RNO_303 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_412, B => memoryro_108, C => 
        memorya412_Z, D => memorya108_Z, Y => memoryror_4);
    
    memoryrff_124 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_124, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_124);
    
    memorya270_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya273_4_Z, B => memorya46_3_Z, Y => 
        memorya270_6_Z);
    
    memoryrff_86_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya86_Z, B => WriteEnable, Y => 
        memorywre_86);
    
    memoryrff_465 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_465, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_465);
    
    memorya6 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya102_1_Z, B => memorya4_6_Z, C => 
        InternalAddr2Memory(8), D => memorya102_3_Z, Y => 
        memorya6_Z);
    
    memorya417 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya353_1_Z, 
        C => memorya353_6_Z, D => memorya498_3_Z, Y => 
        memorya417_Z);
    
    memoryrff_131 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_131, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_131);
    
    memorya67_2 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(2), Y => memorya67_2_Z);
    
    memoryrff_32 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_32, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_32);
    
    memorya270 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya102_1_Z, 
        C => memorya264_1_Z, D => memorya270_6_Z, Y => 
        memorya270_Z);
    
    memorya401 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya369_1_Z, 
        C => memorya336_6_Z, D => memorya498_3_Z, Y => 
        memorya401_Z);
    
    memorya424 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya45_2_Z, C
         => memorya360_6_Z, D => memorya498_3_Z, Y => 
        memorya424_Z);
    
    memorya392 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya393_6_Z, B => memorya370_3_Z, C => 
        InternalAddr2Memory(6), D => memorya395_2_Z, Y => 
        memorya392_Z);
    
    memorya386_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(1), Y => memorya386_1_Z);
    
    memoryrff_391 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_391, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_391);
    
    memory_memory_0_0_sr_RNO_371 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya261_0_Z, B => memorya268_6_Z, C => 
        memorya264_1_Z, Y => memorya269);
    
    memory_memory_0_0_sr_RNO_193 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_207, B => memoryro_399, C => 
        memorya399_Z, D => memorya207_Z, Y => memoryror_131);
    
    memoryrff_157 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_157, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_157);
    
    memoryrff_12_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya68_2_Z, C => 
        memorya12_0_Z, D => memorya4_6_Z, Y => memorywre_12);
    
    memorya308 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya68_2_Z, B => memorya304_4_Z, C => 
        memorya276_0_Z, D => memorya305_2_Z, Y => memorya308_Z);
    
    memorya116 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya116_4_Z, B => memorya116_1_Z, C => 
        memorya20_0_Z, D => memorya116_2_Z, Y => memorya116_Z);
    
    memoryrff_398_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya398_Z, B => WriteEnable, Y => 
        memorywre_398);
    
    memorya315_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya379_1_Z, B => memorya125_2_Z, Y => 
        memorya315_5_Z);
    
    memory_memory_0_0_sr_RNO_382 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya20_6_Z, B => memorya102_1_Z, C => 
        memorya16_0_Z, Y => memorya22);
    
    memory_memory_0_0_sr_RNO_159 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_282, B => memoryro_170, C => 
        memorya282_Z, D => memorya170_Z, Y => memoryror_172);
    
    memoryrff_177 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_177, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_177);
    
    memory_memory_0_0_sr_RNO_150 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_166, B => memoryro_470, C => 
        memorya470_Z, D => memorya166_Z, Y => memoryror_170);
    
    memoryrff_489 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_489, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_489);
    
    memoryrff_268_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya268_Z, B => WriteEnable, Y => 
        memorywre_268);
    
    memoryrff_195 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_195, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_195);
    
    memoryrff_436 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_436, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_436);
    
    memorya499 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(3), B => memorya379_4_Z, 
        C => memorya482_2_Z, D => memorya499_5_Z, Y => 
        memorya499_Z);
    
    memorya393 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya121_1_Z, 
        C => memorya393_6_Z, D => memorya498_3_Z, Y => 
        memorya393_Z);
    
    memorya110 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya84_2_Z, C
         => memorya102_4_Z, D => memorya110_5_Z, Y => 
        memorya110_Z);
    
    memory_memory_0_0_sr_RNO_6 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_433, B => memoryror_435, C => 
        memoryror_432, D => memoryror_434, Y => memoryror_492);
    
    memory_memory_0_0_sr_RNO_116 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_189, B => memoryro_461, C => 
        memorya461_Z, D => memorya189_Z, Y => memoryror_198);
    
    memoryrff_360_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya360_Z, B => WriteEnable, Y => 
        memorywre_360);
    
    memoryrff_353 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_353, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_353);
    
    memorya368_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(2), Y => memorya368_4_Z);
    
    memorya25 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya25_3_Z, B => memorya121_1_Z, C => 
        memorya52_4, D => memorya21_0_Z, Y => memorya25_Z);
    
    memory_memory_0_0_sr_RNO_163 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_172, B => memoryro_364, C => 
        memorya364_Z, D => memorya172_Z, Y => memoryror_164);
    
    memoryrff_373 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_373, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_373);
    
    memoryrff_114_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya114_Z, B => WriteEnable, Y => 
        memorywre_114);
    
    memorya143_0 : CFG3
      generic map(INIT => x"04")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(7), C => InternalAddr2Memory(8), Y
         => memorya143_0_Z);
    
    memory_memory_0_0_sr_RNO_94 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_196, B => memoryro_276, C => 
        memorya276_Z, D => memorya196_Z, Y => memoryror_217);
    
    memoryrff_94 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_94, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_94);
    
    memorya24 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya125_2_Z, B => memorya25_3_Z, C => 
        memorya52_4, D => memorya20_0_Z, Y => memorya24_Z);
    
    memoryrff_44_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya52_2_Z, B => WriteEnable, C => 
        memorya45_6_Z, D => memorya12_0_Z, Y => memorywre_44);
    
    memoryrff_109 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_109, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_109);
    
    memorya90 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya362_1_Z, B => memorya86_2_Z, C => 
        memorya68_4_Z, D => memorya10_0_Z, Y => memorya90_Z);
    
    memoryrff_226 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_226, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_226);
    
    memorya359 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya68_3_Z, C
         => memorya368_2_Z, D => memorya487_5_Z, Y => 
        memorya359_Z);
    
    memorya370_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(1), Y => memorya370_1_Z);
    
    memorya280 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya280_6_Z, B => memorya280_0_Z, C => 
        memorya370_3_Z, Y => memorya280_Z);
    
    memoryrff_369_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya369_Z, B => WriteEnable, Y => 
        memorywre_369);
    
    memorya349 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya29_3_Z, C
         => memorya368_2_Z, D => memorya381_5_Z, Y => 
        memorya349_Z);
    
    memory_memory_0_0_sr_RNO_338 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_278, B => memoryro_22, C => 
        memorya278_Z, D => memorya22, Y => memoryror_26);
    
    memoryrff_228_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya228_Z, B => WriteEnable, Y => 
        memorywre_228);
    
    memoryrff_111_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya463_5_Z, B => memorya111_0_Z, C => 
        WriteEnable, D => memorya102_4_Z, Y => memorywre_111);
    
    memorya45_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(1), Y => memorya45_3_Z);
    
    memoryrff_168 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_168, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_168);
    
    memorya273_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya273_4_Z, B => memorya368_4_Z, Y => 
        memorya273_6_Z);
    
    memory_memory_0_0_sr_RNO_34 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_245, B => memoryror_247, C => 
        memoryror_244, D => memoryror_246, Y => memoryror_445);
    
    memory_memory_0_0_sr_RNO_142 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_316, B => memoryro_252, C => 
        memorya316_Z, D => memorya252_Z, Y => memoryror_244);
    
    memoryrff_478_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya478_Z, B => WriteEnable, Y => 
        memorywre_478);
    
    memoryrff_320_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya320_Z, B => WriteEnable, Y => 
        memorywre_320);
    
    memoryrff_267 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_267, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_267);
    
    memoryrff_215_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya215_Z, B => WriteEnable, Y => 
        memorywre_215);
    
    memoryrff_115_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya115_Z, B => WriteEnable, Y => 
        memorywre_115);
    
    memoryrff_9_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya57_3_Z, C => 
        memorya9_0_Z, D => memorya4_6_Z, Y => memorywre_9);
    
    memoryrff_78_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya78_Z, B => WriteEnable, Y => 
        memorywre_78);
    
    memoryrff_310 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_310, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_310);
    
    memoryrff_248 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_248, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_248);
    
    memory_memory_0_0_sr_RNO_118 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_220, B => memoryro_268, C => 
        memorya268_Z, D => memorya220_Z, Y => memoryror_196);
    
    memoryrff_271_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya271_Z, B => WriteEnable, Y => 
        memorywre_271);
    
    memoryrff_212_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya212_Z, B => WriteEnable, Y => 
        memorywre_212);
    
    memoryrff_85_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya85_Z, B => WriteEnable, Y => 
        memorywre_85);
    
    memoryrff_329_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya329_Z, B => WriteEnable, Y => 
        memorywre_329);
    
    memory_memory_0_0_sr_RNO_351 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya20_6_Z, B => memorya370_1_Z, C => 
        memorya10_0_Z, Y => memorya18);
    
    memoryrff_493 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_493, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_493);
    
    memoryrff_490 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_490, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_490);
    
    memorya68_2 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(1), Y => memorya68_2_Z);
    
    memoryrff_460_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya460_Z, B => WriteEnable, Y => 
        memorywre_460);
    
    memorya329 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya121_1_Z, 
        C => memorya368_2_Z, D => memorya393_6_Z, Y => 
        memorya329_Z);
    
    memoryrff_77_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya77_Z, B => WriteEnable, Y => 
        memorywre_77);
    
    memoryrff_206_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya206_Z, B => WriteEnable, Y => 
        memorywre_206);
    
    memoryrff_373_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya373_Z, B => WriteEnable, Y => 
        memorywre_373);
    
    memory_memory_0_0_sr_RNO_9 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_423, B => memoryror_421, C => 
        memoryror_422, D => memoryror_420, Y => memoryror_489);
    
    memoryrff_162_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya162_Z, B => WriteEnable, Y => 
        memorywre_162);
    
    \memory_memory_0_0_OLDA_RNICPU31[25]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(25), C => 
        memory_memory_0_0_OLDA_Z(25), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(25));
    
    memoryrff_69 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_69, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_69);
    
    memory_memory_0_0_sr_RNO_300 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_269, B => memoryro_61, C => 
        memorya269, D => memorya61_Z, Y => memoryror_6);
    
    memory_memory_0_0_sr_RNO_297 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_6, B => memoryro_262, C => 
        memorya262_Z, D => memorya6_Z, Y => memoryror_10);
    
    memoryrff_435 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_435, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_435);
    
    memoryrff_194 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_194, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_194);
    
    memoryrff_254_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya254_Z, B => WriteEnable, Y => 
        memorywre_254);
    
    memoryrff_234_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya234_Z, B => WriteEnable, Y => 
        memorywre_234);
    
    memorya208 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya86_2_Z, C
         => memorya162_2_Z, D => memorya336_6_Z, Y => 
        memorya208_Z);
    
    memorya501 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(3), B => memorya369_3_Z, 
        C => memorya373_5_Z, D => memorya482_2_Z, Y => 
        memorya501_Z);
    
    memoryrff_409 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_409, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_409);
    
    memory_memory_0_0_sr_RNO_3 : CFG4
      generic map(INIT => x"FFFB")

      port map(A => memoryror_483, B => memoryror_504_1, C => 
        memoryror_482, D => memoryror_481, Y => memoryror_504);
    
    memorya202 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya362_1_Z, 
        C => memorya202_6_Z, D => memorya482_2_Z, Y => 
        memorya202_Z);
    
    memoryrff_420_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya420_Z, B => WriteEnable, Y => 
        memorywre_420);
    
    memoryrff_121 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_121, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_121);
    
    memory_memory_0_0_sr_RNO_72 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_14, B => memoryror_13, C => 
        memoryror_12, D => memoryror_15, Y => memoryror_387);
    
    memory_memory_0_0_sr_RNO_267 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_375, B => memoryro_119, C => 
        memorya375_Z, D => memorya119, Y => memoryror_126);
    
    memorya451 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_1_Z, B => InternalAddr2Memory(5), 
        C => memorya355_6_Z, D => memorya482_2_Z, Y => 
        memorya451_Z);
    
    memoryrff_39 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_39, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_39);
    
    memoryrff_351 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_351, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_351);
    
    memoryrff_122_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya122_Z, B => WriteEnable, Y => 
        memorywre_122);
    
    memorya211_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya20_3_Z, B => InternalAddr2Memory(8), Y
         => memorya211_0_Z);
    
    memorya441 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya54_2_Z, B => memorya441_6_Z, C => 
        InternalAddr2Memory(6), D => memorya121_1_Z, Y => 
        memorya441_Z);
    
    memorya358_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya370_3_Z, B => memorya68_3_Z, Y => 
        memorya358_6_Z);
    
    memorya358 : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory(7), B => memorya102_5_Z, 
        C => memorya358_6_Z, Y => memorya358_Z);
    
    memoryrff_178_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya178_Z, B => WriteEnable, Y => 
        memorywre_178);
    
    memory_memory_0_0_sr_RNO_289 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_309, B => memoryro_53, C => 
        memorya309_Z, D => memorya53_Z, Y => memoryror_59);
    
    memory_memory_0_0_sr_RNO_285 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_318, B => memoryro_190, C => 
        memorya318_Z, D => memorya190_Z, Y => memoryror_55);
    
    memoryrff_371 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_371, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_371);
    
    memorya348 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya29_3_Z, B => InternalAddr2Memory(7), C
         => memorya348_5_Z, D => memorya370_3_Z, Y => 
        memorya348_Z);
    
    memoryrff_155 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_155, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_155);
    
    memory_memory_0_0_sr_RNO_134 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_306, B => memoryro_114, C => 
        memorya306_Z, D => memorya114_Z, Y => memoryror_240);
    
    memorya4 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya4_0_Z, B => InternalAddr2Memory(8), C
         => memorya84_3_Z, D => memorya4_6_Z, Y => memorya4_Z);
    
    memorya21_0 : CFG3
      generic map(INIT => x"04")

      port map(A => InternalAddr2Memory(1), B => 
        InternalAddr2Memory(4), C => InternalAddr2Memory(8), Y
         => memorya21_0_Z);
    
    memoryrff_426 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_426, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_426);
    
    memoryrff_175 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_175, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_175);
    
    memorya149_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya403_2_Z, B => memorya117_1_Z, Y => 
        memorya149_5_Z);
    
    memory_memory_0_0_sr_RNO_248 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_102, B => memoryro_358, C => 
        memorya358_Z, D => memorya102_Z, Y => memoryror_106);
    
    memoryrff_287_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya287_Z, B => WriteEnable, Y => 
        memorywre_287);
    
    memory_memory_0_0_sr_RNO_11 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_429, B => memoryror_431, C => 
        memoryror_428, D => memoryror_430, Y => memoryror_491);
    
    memory_memory_0_0_sr_RNO_272 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_374, B => memoryro_118, C => 
        memorya374_Z, D => memorya118_Z, Y => memoryror_122);
    
    memoryrff_147 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_147, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_147);
    
    memorya273 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya369_1_Z, B => InternalAddr2Memory(7), 
        C => memorya273_6_Z, D => memorya369_3_Z, Y => 
        memorya273_Z);
    
    memoryrff_140_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya140_Z, B => WriteEnable, Y => 
        memorywre_140);
    
    memoryrff_46_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya46_Z, B => WriteEnable, Y => 
        memorywre_46);
    
    memorya95 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya86_2_Z, C
         => memorya68_4_Z, D => memorya463_5_Z, Y => memorya95_Z);
    
    memorya116_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(3), Y => memorya116_4_Z);
    
    memorya421 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya117_1_Z, B => InternalAddr2Memory(6), 
        C => memorya421_6_Z, D => memorya434_2_Z, Y => 
        memorya421_Z);
    
    memoryrff_138 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_138, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_138);
    
    memorya94 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya84_2_Z, C
         => memorya68_4_Z, D => memorya126_5_Z, Y => memorya94_Z);
    
    memorya487_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya379_1_Z, B => memorya36_1_Z, Y => 
        memorya487_5_Z);
    
    memoryrff_364 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_364, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_364);
    
    memoryrff_296 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_296, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_296);
    
    memorya328 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya77_2_Z, B => InternalAddr2Memory(7), C
         => memorya370_3_Z, D => memorya393_6_Z, Y => 
        memorya328_Z);
    
    memoryrff_463_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya463_Z, B => WriteEnable, Y => 
        memorywre_463);
    
    memoryrff_343 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_343, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_343);
    
    memoryrff_237 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_237, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_237);
    
    memorya316_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(1), Y => memorya316_4_Z);
    
    \memory_memory_0_0_OLDA_RNIERU31[27]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(27), C => 
        memory_memory_0_0_OLDA_Z(27), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(27));
    
    memoryrff_454_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya454_Z, B => WriteEnable, Y => 
        memorywre_454);
    
    memoryrff_106_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya106_Z, B => WriteEnable, Y => 
        memorywre_106);
    
    memory_memory_0_0_sr_RNO_226 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_433, B => memoryro_17, C => 
        memorya433_Z, D => memorya17_Z, Y => memoryror_81);
    
    memoryrff_434_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya434_Z, B => WriteEnable, Y => 
        memorywre_434);
    
    memoryrff_183_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya183_Z, B => WriteEnable, Y => 
        memorywre_183);
    
    memory_memory_0_0_sr_RNO_308 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_174, B => memoryro_302, C => 
        memorya302_Z, D => memorya174_Z, Y => memoryror_39);
    
    memoryrff_449_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya449_Z, B => WriteEnable, Y => 
        memorywre_449);
    
    memorya342_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya370_3_Z, B => memorya20_3_Z, Y => 
        memorya342_6_Z);
    
    memoryrff_385_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya385_Z, B => WriteEnable, Y => 
        memorywre_385);
    
    \memory_memory_0_0_OLDA_RNITUUT[8]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(8), C => 
        memory_memory_0_0_OLDA_Z(8), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(8));
    
    memoryrff_476_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya476_Z, B => WriteEnable, Y => 
        memorywre_476);
    
    memoryrff_453 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_453, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_453);
    
    memoryrff_450 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_450, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_450);
    
    memorya283 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya273_4_Z, B => InternalAddr2Memory(7), 
        C => memorya315_5_Z, D => memorya379_4_Z, Y => 
        memorya283_Z);
    
    memorya260_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(2), Y => memorya260_1_Z);
    
    memorya92 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya364_1_Z, B => memorya86_2_Z, C => 
        memorya68_4_Z, D => memorya20_0_Z, Y => memorya92_Z);
    
    memorya395 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya4_3_Z, C
         => memorya379_4_Z, D => memorya395_5_Z, Y => 
        memorya395_Z);
    
    memoryrff_372_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya372_Z, B => WriteEnable, Y => 
        memorywre_372);
    
    memorya354_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya68_3_Z, B => memorya354_3_Z, Y => 
        memorya354_6_Z);
    
    memorya114 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya370_1_Z, B => memorya116_4_Z, C => 
        memorya116_2_Z, D => memorya10_0_Z, Y => memorya114_Z);
    
    memory_memory_0_0_sr_RNO_347 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya36_6_Z, B => memorya354_1_Z, C => 
        memorya10_0_Z, Y => memorya34);
    
    memoryrff_423_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya423_Z, B => WriteEnable, Y => 
        memorywre_423);
    
    memoryrff_473 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_473, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_473);
    
    memoryrff_470 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_470, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_470);
    
    \memory_memory_0_0_OLDA_RNISTUT[7]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(7), C => 
        memory_memory_0_0_OLDA_Z(7), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(7));
    
    memorya258_0 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(1), Y => memorya258_0_Z);
    
    memoryrff_65 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_65, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_65);
    
    memoryrff_216_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya216_Z, B => WriteEnable, Y => 
        memorywre_216);
    
    memorya56_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya125_2_Z, B => InternalAddr2Memory(8), 
        Y => memorya56_0_Z);
    
    memorya395_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(3), Y => memorya395_2_Z);
    
    memorya368_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya68_2_Z, B => memorya368_4_Z, Y => 
        memorya368_6_Z);
    
    memory_memory_0_0_sr_RNO_243 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_417, B => memoryro_1, C => 
        memorya417_Z, D => memorya1_Z, Y => memoryror_65);
    
    memoryrff_67 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_67, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_67);
    
    memoryrff_190_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya190_Z, B => WriteEnable, Y => 
        memorywre_190);
    
    memoryrff_154 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_154, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_154);
    
    memoryrff_149_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya149_Z, B => WriteEnable, Y => 
        memorywre_149);
    
    memoryrff_425 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_425, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_425);
    
    memory_memory_0_0_sr_RNO_252 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_400, B => memoryro_208, C => 
        memorya400_Z, D => memorya208_Z, Y => memoryror_98);
    
    memorya1_0 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(1), Y => memorya1_0_Z);
    
    memoryrff_174 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_174, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_174);
    
    memorya258 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya258_0_Z, B => memorya257_6_Z, C => 
        InternalAddr2Memory(7), D => memorya354_3_Z, Y => 
        memorya258_Z);
    
    memory_memory_0_0_sr_RNO_59 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_66, B => memoryror_64, C => 
        memoryror_67, D => memoryror_65, Y => memoryror_400);
    
    memorya252 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya68_2_Z, C
         => memorya380_5_Z, D => memorya482_2_Z, Y => 
        memorya252_Z);
    
    memorya248 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya116_2_Z, B => memorya128_0_Z, C => 
        memorya125_2_Z, Y => memorya248_Z);
    
    memoryrff_81_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya81_Z, B => WriteEnable, Y => 
        memorywre_81);
    
    memorya20_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya68_2_Z, B => InternalAddr2Memory(8), Y
         => memorya20_0_Z);
    
    memory_memory_0_0_sr_RNO_119 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_475, B => memoryro_27, C => 
        memorya475_Z, D => memorya27_Z, Y => memoryror_197);
    
    memorya509 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya116_2_Z, B => InternalAddr2Memory(1), 
        C => memorya381_5_Z, D => memorya498_3_Z, Y => 
        memorya509_Z);
    
    memory_memory_0_0_sr_RNO_110 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_233, B => memoryro_489, C => 
        memorya489_Z, D => memorya233_Z, Y => memoryror_237);
    
    memorya242 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya116_2_Z, B => memorya370_1_Z, C => 
        memorya162_2_Z, D => memorya3_0_Z, Y => memorya242_Z);
    
    memoryrff_35 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_35, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_35);
    
    memorya19 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya19_0_Z, B => InternalAddr2Memory(8), C
         => memorya379_1_Z, D => memorya20_6_Z, Y => memorya19_Z);
    
    memoryrff_191 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_191, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_191);
    
    memoryrff_18_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya370_1_Z, B => WriteEnable, C => 
        memorya20_6_Z, D => memorya10_0_Z, Y => memorywre_18);
    
    memoryrff_499_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya499_Z, B => WriteEnable, Y => 
        memorywre_499);
    
    memoryrff_37 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_37, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_37);
    
    memorya414 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya30_3_Z, B => InternalAddr2Memory(6), C
         => memorya126_5_Z, D => memorya498_3_Z, Y => 
        memorya414_Z);
    
    memoryrff_78 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_78, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_78);
    
    memoryrff_45_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya45_Z, B => WriteEnable, Y => 
        memorywre_45);
    
    memorya211_3 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(2), Y => memorya211_3_Z);
    
    memoryrff_401_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya401_Z, B => WriteEnable, Y => 
        memorywre_401);
    
    memory_memory_0_0_sr_RNO_56 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_71, B => memoryror_69, C => 
        memoryror_70, D => memoryror_68, Y => memoryror_401);
    
    memoryrff_17_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya17_Z, B => WriteEnable, Y => 
        memorywre_17);
    
    memoryrff_505 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_505, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_505);
    
    memoryrff_11 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_11, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_11);
    
    memory_memory_0_0_sr_RNO_89 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_159, B => memoryro_479, C => 
        memorya479_Z, D => memorya159_Z, Y => memoryror_211);
    
    memoryrff_160 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_160, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_160);
    
    memoryrff_496 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_496, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_496);
    
    memory_memory_0_0_sr_RNO_62 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_98, B => memoryror_96, C => 
        memoryror_99, D => memoryror_97, Y => memoryror_408);
    
    memory_memory_0_0_sr_RNO_183 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_502, B => memoryro_134, C => 
        memorya502_Z, D => memorya134_Z, Y => memoryror_138);
    
    memory_memory_0_0_sr_RNO_104 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_157, B => memoryro_493, C => 
        memorya493_Z, D => memorya157_Z, Y => memoryror_230);
    
    memoryrff_341 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_341, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_341);
    
    memoryrff_283 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_283, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_283);
    
    memorya228 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya36_1_Z, C
         => memorya356_6_Z, D => memorya482_2_Z, Y => 
        memorya228_Z);
    
    memorya266_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya362_1_Z, B => InternalAddr2Memory(7), 
        Y => memorya266_0_Z);
    
    memorya117_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(2), Y => memorya117_1_Z);
    
    memory_memory_0_0_sr_RNO_274 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_116, B => memoryro_500, C => 
        memorya500_Z, D => memorya116_Z, Y => memoryror_121);
    
    memorya356_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya68_2_Z, B => memorya68_3_Z, Y => 
        memorya356_6_Z);
    
    memorya222 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya30_3_Z, C
         => memorya126_5_Z, D => memorya482_2_Z, Y => 
        memorya222_Z);
    
    memoryrff_468_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya468_Z, B => WriteEnable, Y => 
        memorywre_468);
    
    memoryrff_334 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_334, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_334);
    
    memorya290 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya354_1_Z, B => InternalAddr2Memory(7), 
        C => memorya289_6_Z, D => memorya370_3_Z, Y => 
        memorya290_Z);
    
    memoryrff_511 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_511, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_511);
    
    memory_memory_0_0_sr_RNO_23 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_214, B => memoryror_215, C => 
        memoryror_212, D => memoryror_213, Y => memoryror_437);
    
    memoryrff_154_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya154_Z, B => WriteEnable, Y => 
        memorywre_154);
    
    memoryrff_145 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_145, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_145);
    
    memorya233_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya41_3_Z, B => InternalAddr2Memory(8), Y
         => memorya233_0_Z);
    
    memoryrff_315 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_315, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_315);
    
    memoryrff_199_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya199_0_Z, B => memorya455_5_Z, C => 
        WriteEnable, D => memorya167_3_Z, Y => memorywre_199);
    
    memoryrff_134_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya134_Z, B => WriteEnable, Y => 
        memorywre_134);
    
    memorya274 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya370_1_Z, B => InternalAddr2Memory(7), 
        C => memorya273_6_Z, D => memorya370_3_Z, Y => 
        memorya274_Z);
    
    memoryrff_256 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_256, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_256);
    
    memoryrff_128 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_128, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_128);
    
    memoryrff_371_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya371_Z, B => WriteEnable, Y => 
        memorywre_371);
    
    memorya393_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya4_3_Z, B => memorya57_3_Z, Y => 
        memorya393_6_Z);
    
    memory_memory_0_0_sr_RNO_86 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_330, B => memoryro_218, C => 
        memorya330_Z, D => memorya218_Z, Y => memoryror_220);
    
    memorya369_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(0), Y => memorya369_1_Z);
    
    memory_memory_0_0_sr_RNO_363 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya68_2_Z, B => memorya12_0_Z, C => 
        memorya4_6_Z, Y => memorya12);
    
    memoryrff_261_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya261_Z, B => WriteEnable, Y => 
        memorywre_261);
    
    memory_memory_0_0_sr_RNO_175 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_150, B => memoryro_486, C => 
        memorya486_Z, D => memorya150_Z, Y => memoryror_154);
    
    memoryrff_276 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_276, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_276);
    
    memorya364_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya370_3_Z, B => memorya45_3_Z, Y => 
        memorya364_6_Z);
    
    memoryrff_227 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_227, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_227);
    
    memorya30 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya30_3_Z, C
         => memorya52_4, D => memorya126_5_Z, Y => memorya30_Z);
    
    memory_memory_0_0_sr_RNO_375 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya292_6_Z, B => memorya305_2_Z, C => 
        memorya261_0_Z, Y => memorya293);
    
    memory_memory_0_0_sr_RNO_271 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_127, B => memoryro_383, C => 
        memorya383_Z, D => memorya127_Z, Y => memoryror_115);
    
    memoryrff_319 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_319, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_319);
    
    memoryrff_151_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya151_Z, B => WriteEnable, Y => 
        memorywre_151);
    
    memorya268_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya364_1_Z, B => InternalAddr2Memory(7), 
        Y => memorya268_0_Z);
    
    memorya13_0 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(1), Y => memorya13_0_Z);
    
    memoryrff_131_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya131_Z, B => WriteEnable, Y => 
        memorywre_131);
    
    memory_memory_0_0_sr_RNO_311 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_76, B => memoryro_428, C => 
        memorya428_Z, D => memorya76_Z, Y => memoryror_36);
    
    \memory_memory_0_0_OLDA_RNIFRT31[19]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(19), C => 
        memory_memory_0_0_OLDA_Z(19), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(19));
    
    \memory_memory_0_0_OLDA_RNIBOU31[24]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(24), C => 
        memory_memory_0_0_OLDA_Z(24), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(24));
    
    \memory_memory_0_0_OLDA_RNIANU31[23]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(23), C => 
        memory_memory_0_0_OLDA_Z(23), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(23));
    
    memoryrff_363_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya363_Z, B => WriteEnable, Y => 
        memorywre_363);
    
    memoryrff_116_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya116_Z, B => WriteEnable, Y => 
        memorywre_116);
    
    memorya264_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(3), Y => memorya264_1_Z);
    
    memoryrff_81 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_81, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_81);
    
    memoryrff_428_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya428_Z, B => WriteEnable, Y => 
        memorywre_428);
    
    memoryrff_255_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya255_Z, B => WriteEnable, Y => 
        memorywre_255);
    
    memoryrff_2 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_2, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_2);
    
    memorya475 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_4_Z, B => InternalAddr2Memory(5), 
        C => memorya315_5_Z, D => memorya482_2_Z, Y => 
        memorya475_Z);
    
    memory_memory_0_0_sr_RNO_270 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_385, B => memoryro_49, C => 
        memorya385_Z, D => memorya49_Z, Y => memoryror_113);
    
    memoryrff_235_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya235_Z, B => WriteEnable, Y => 
        memorywre_235);
    
    memoryrff_155_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya155_Z, B => WriteEnable, Y => 
        memorywre_155);
    
    memorya370_3 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(0), Y => memorya370_3_Z);
    
    \memory_memory_0_0_OLDA[18]\ : SLE
      port map(D => \InternalDataFromMem\(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(18));
    
    memoryrff_135_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya135_Z, B => WriteEnable, Y => 
        memorywre_135);
    
    memorya16_0 : CFG3
      generic map(INIT => x"04")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(4), C => InternalAddr2Memory(8), Y
         => memorya16_0_Z);
    
    memoryrff_252_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya252_Z, B => WriteEnable, Y => 
        memorywre_252);
    
    memoryrff_221_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya221_Z, B => WriteEnable, Y => 
        memorywre_221);
    
    memoryrff_232_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya232_Z, B => WriteEnable, Y => 
        memorywre_232);
    
    memorya31_0 : CFG2
      generic map(INIT => x"4")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(4), Y => memorya31_0_Z);
    
    memorya319 : CFG4
      generic map(INIT => x"8000")

      port map(A => InternalAddr2Memory(8), B => memorya54_2_Z, C
         => memorya52_4, D => memorya463_5_Z, Y => memorya319_Z);
    
    memorya284 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya273_4_Z, B => memorya68_2_Z, C => 
        memorya268_0_Z, D => memorya278_2_Z, Y => memorya284_Z);
    
    memoryrff_509_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya509_Z, B => WriteEnable, Y => 
        memorywre_509);
    
    memoryrff_307_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya307_Z, B => WriteEnable, Y => 
        memorywre_307);
    
    memory_memory_0_0_sr_RNO_92 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_211, B => memoryro_339, C => 
        memorya339_Z, D => memorya211_Z, Y => memoryror_216);
    
    memoryrff_384_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya384_Z, B => WriteEnable, Y => 
        memorywre_384);
    
    \memory_memory_0_0_OLDA_RNIPQUT[4]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(4), C => 
        memory_memory_0_0_OLDA_Z(4), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(4));
    
    memoryrff_323_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya323_Z, B => WriteEnable, Y => 
        memorywre_323);
    
    memoryrff_443 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_443, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_443);
    
    memoryrff_440 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_440, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_440);
    
    memoryrff_70 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_70, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_70);
    
    memory_memory_0_0_sr_RNO_254 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_367, B => memoryro_111, C => 
        memorya367_Z, D => memorya111, Y => memoryror_99);
    
    memoryrff_495 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_495, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_495);
    
    memoryrff_168_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya168_Z, B => WriteEnable, Y => 
        memorywre_168);
    
    memorya319_0 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(6), Y => memorya52_4);
    
    memory_memory_0_0_sr_RNO_287 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_444, B => memoryro_92, C => 
        memorya444_Z, D => memorya92_Z, Y => memoryror_52);
    
    memoryrff_64 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_64, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_64);
    
    memorya485 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya84_3_Z, B => InternalAddr2Memory(4), C
         => memorya101_5_Z, D => memorya498_3_Z, Y => 
        memorya485_Z);
    
    memory_memory_0_0_sr_RNO_32 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_241, B => memoryror_242, C => 
        memoryror_240, D => memoryror_243, Y => memoryror_444);
    
    memory_memory_0_0_sr_RNO_122 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_328, B => memoryro_184, C => 
        memorya328_Z, D => memorya184_Z, Y => memoryror_207);
    
    memoryrff_99_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya99_Z, B => WriteEnable, Y => 
        memorywre_99);
    
    memoryrff_39_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya39_Z, B => WriteEnable, Y => 
        memorywre_39);
    
    memorya402 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya370_1_Z, 
        C => memorya338_6_Z, D => memorya498_3_Z, Y => 
        memorya402_Z);
    
    memory_memory_0_0_sr_RNO_44 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_137, B => memoryror_139, C => 
        memoryror_136, D => memoryror_138, Y => memoryror_418);
    
    memoryrff_151 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_151, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_151);
    
    memoryrff_203 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_203, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_203);
    
    memory_memory_0_0_sr_RNO_155 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_322, B => memoryro_34, C => 
        memorya322_Z, D => memorya34, Y => memoryror_160);
    
    memoryrff_144 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_144, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_144);
    
    \memory_memory_0_0_OLDA_RNIEQT31[18]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(18), C => 
        memory_memory_0_0_OLDA_Z(18), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(18));
    
    memory_memory_0_0_sr_RNO_355 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya51_6_Z, B => memorya54_2_Z, C => 
        memorya20_0_Z, Y => memorya48);
    
    memoryrff_171 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_171, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_171);
    
    memory_memory_0_0_sr_RNO_251 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_357, B => memoryro_101, C => 
        memorya357_Z, D => memorya101_Z, Y => memoryror_107);
    
    memoryrff_130 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_130, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_130);
    
    memorya464_0 : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory(5), B => memorya86_2_Z, C
         => memorya498_3_Z, Y => memorya464_0_Z);
    
    memorya460 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya364_1_Z, B => InternalAddr2Memory(5), 
        C => memorya364_6_Z, D => memorya482_2_Z, Y => 
        memorya460_Z);
    
    memory_memory_0_0_sr_RNO_177 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_415, B => memoryro_223, C => 
        memorya415_Z, D => memorya223_Z, Y => memoryror_147);
    
    memoryrff_128_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya68_3_Z, C => 
        memorya273_4_Z, D => memorya128_0_Z, Y => memorywre_128);
    
    memoryrff_411_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya411_Z, B => WriteEnable, Y => 
        memorywre_411);
    
    memoryrff_407_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya407_Z, B => WriteEnable, Y => 
        memorywre_407);
    
    memorya430 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya46_3_Z, C
         => memorya110_5_Z, D => memorya498_3_Z, Y => 
        memorya430_Z);
    
    memorya42_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya362_1_Z, B => InternalAddr2Memory(8), 
        Y => memorya42_0_Z);
    
    memory_memory_0_0_sr_RNO_250 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_403, B => memoryro_99, C => 
        memorya403_Z, D => memorya99_Z, Y => memoryror_104);
    
    memoryrff_456 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_456, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_456);
    
    memoryrff_34 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_34, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_34);
    
    memorya306 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya305_2_Z, B => memorya306_6_Z, C => 
        InternalAddr2Memory(7), D => memorya370_1_Z, Y => 
        memorya306_Z);
    
    memoryrff_4 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_4, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_4);
    
    memorya70 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya84_2_Z, B => memorya68_6_Z, C => 
        InternalAddr2Memory(8), D => memorya102_1_Z, Y => 
        memorya70_Z);
    
    memoryrff_476 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_476, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_476);
    
    memorya474_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya86_2_Z, B => memorya362_1_Z, Y => 
        memorya474_5_Z);
    
    memorya199_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya4_3_Z, B => InternalAddr2Memory(8), Y
         => memorya199_0_Z);
    
    memoryrff_92_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya92_Z, B => WriteEnable, Y => 
        memorywre_92);
    
    memoryrff_32_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya32_Z, B => WriteEnable, Y => 
        memorywre_32);
    
    memoryrff_324 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_324, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_324);
    
    memorya411 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya25_3_Z, B => InternalAddr2Memory(6), C
         => memorya315_5_Z, D => memorya498_3_Z, Y => 
        memorya411_Z);
    
    memorya205 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya77_2_Z, B => memorya117_1_Z, C => 
        memorya199_0_Z, D => memorya193_2_Z, Y => memorya205_Z);
    
    memory_memory_0_0_sr_RNO_360 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya432_0_Z, B => memorya368_6_Z, Y => 
        memorya432);
    
    memoryrff_41_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya41_Z, B => WriteEnable, Y => 
        memorywre_41);
    
    memoryrff_198 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_198, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_198);
    
    memory_memory_0_0_sr_RNO_20 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_222, B => memoryror_221, C => 
        memoryror_220, D => memoryror_223, Y => memoryror_439);
    
    memoryrff_466_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya466_Z, B => WriteEnable, Y => 
        memorywre_466);
    
    memoryrff_0 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_0, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_0);
    
    memorya318 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya305_2_Z, B => memorya126_5_Z, C => 
        InternalAddr2Memory(7), D => memorya318_4_Z, Y => 
        memorya318_Z);
    
    memory_memory_0_0_sr_RNO_4 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_439, B => memoryror_436, C => 
        memoryror_438, D => memoryror_437, Y => memoryror_493);
    
    memoryrff_362_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya362_Z, B => WriteEnable, Y => 
        memorywre_362);
    
    memoryrff_308_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya308_Z, B => WriteEnable, Y => 
        memorywre_308);
    
    memoryrff_297 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_297, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_297);
    
    memorya463_4 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(4), Y => memorya463_4_Z);
    
    memorya498_3 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(7), Y => memorya498_3_Z);
    
    memoryrff_274_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya274_Z, B => WriteEnable, Y => 
        memorywre_274);
    
    memoryrff_445_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya445_Z, B => WriteEnable, Y => 
        memorywre_445);
    
    memoryrff_246 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_246, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_246);
    
    memorya103 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya87_0, B => memorya102_4_Z, C => 
        memorya487_5_Z, Y => memorya103_Z);
    
    memory_memory_0_0_sr_RNO_349 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya298_6_Z, B => memorya305_2_Z, C => 
        memorya266_0_Z, Y => memorya298);
    
    memory_memory_0_0_sr_RNO_228 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_206, B => memoryro_334, C => 
        memorya334_Z, D => memorya206_Z, Y => memoryror_71);
    
    memory_memory_0_0_sr_RNO_212 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_327, B => memoryro_71, C => 
        memorya327_Z, D => memorya71_Z, Y => memoryror_94);
    
    memoryrff_426_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya426_Z, B => WriteEnable, Y => 
        memorywre_426);
    
    memoryrff_187_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya187_Z, B => WriteEnable, Y => 
        memorywre_187);
    
    memorya91 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya67_2_Z, C
         => memorya68_4_Z, D => memorya315_5_Z, Y => memorya91_Z);
    
    memory_memory_0_0_sr_RNO_157 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_153, B => memoryro_441, C => 
        memorya441_Z, D => memorya153_Z, Y => memoryror_173);
    
    memoryrff_322_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya322_Z, B => WriteEnable, Y => 
        memorywre_322);
    
    memoryrff_461 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_461, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_461);
    
    memorya32 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya52_2_Z, B => InternalAddr2Memory(8), C
         => memorya36_6_Z, D => memorya57_3_Z, Y => memorya32_Z);
    
    memory_memory_0_0_sr_RNO_344 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya368_0_Z, B => memorya368_6_Z, Y => 
        memorya368);
    
    memoryrff_317_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya317_Z, B => WriteEnable, Y => 
        memorywre_317);
    
    memoryrff_256_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya256_Z, B => WriteEnable, Y => 
        memorywre_256);
    
    memoryrff_236_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya236_Z, B => WriteEnable, Y => 
        memorywre_236);
    
    memoryrff_261 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_261, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_261);
    
    memoryrff_23_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya23_Z, B => WriteEnable, Y => 
        memorywre_23);
    
    memoryrff_455 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_455, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_455);
    
    memorya171 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya289_4_Z, 
        C => memorya211_3_Z, D => memorya299_5_Z, Y => 
        memorya171_Z);
    
    memoryrff_289_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya289_Z, B => WriteEnable, Y => 
        memorywre_289);
    
    memory_memory_0_0_sr_RNO_346 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya20_6_Z, B => memorya57_3_Z, C => 
        memorya16_0_Z, Y => memorya16);
    
    memoryrff_475 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_475, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_475);
    
    memorya452 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya68_1_Z, C
         => memorya356_6_Z, D => memorya498_3_Z, Y => 
        memorya452_Z);
    
    memoryrff_282 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_282, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_282);
    
    memorya442 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya54_2_Z, B => memorya498_6_Z, C => 
        InternalAddr2Memory(6), D => memorya362_1_Z, Y => 
        memorya442_Z);
    
    memory_memory_0_0_sr_RNO_171 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_237, B => memoryro_397, C => 
        memorya397_Z, D => memorya237_Z, Y => memoryror_150);
    
    memoryrff_210 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_210, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_210);
    
    memory_memory_0_0_sr_RNO_58 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_77, B => memoryror_79, C => 
        memoryror_76, D => memoryror_78, Y => memoryror_403);
    
    memoryrff_495_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya495_Z, B => WriteEnable, Y => 
        memorywre_495);
    
    memorya370 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya370_1_Z, 
        C => memorya116_2_Z, D => memorya370_6_Z, Y => 
        memorya370_Z);
    
    memoryrff_120 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_120, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_120);
    
    memory_memory_0_0_sr_RNO_368 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya57_3_Z, B => memorya9_0_Z, C => 
        memorya4_6_Z, Y => memorya9);
    
    memorya261_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya117_1_Z, B => InternalAddr2Memory(7), 
        Y => memorya261_0_Z);
    
    memory_memory_0_0_sr_RNO_327 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_146, B => memoryro_466, C => 
        memorya466_Z, D => memorya146_Z, Y => memoryror_16);
    
    memoryrff_474_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya474_Z, B => WriteEnable, Y => 
        memorywre_474);
    
    memorya372_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya370_3_Z, B => memorya84_3_Z, Y => 
        memorya372_6_Z);
    
    memoryrff_361_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya361_Z, B => WriteEnable, Y => 
        memorywre_361);
    
    memoryrff_53_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya53_Z, B => WriteEnable, Y => 
        memorywre_53);
    
    memoryrff_141 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_141, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_141);
    
    memorya356 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya36_1_Z, C
         => memorya356_6_Z, D => memorya368_2_Z, Y => 
        memorya356_Z);
    
    memoryrff_417_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya417_Z, B => WriteEnable, Y => 
        memorywre_417);
    
    memorya75 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya41_3_Z, C
         => memorya68_4_Z, D => memorya331_5_Z, Y => memorya75_Z);
    
    memorya181 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya304_4_Z, 
        C => memorya193_2_Z, D => memorya373_5_Z, Y => 
        memorya181_Z);
    
    memorya346 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya25_3_Z, C
         => memorya370_3_Z, D => memorya474_5_Z, Y => 
        memorya346_Z);
    
    memorya289_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(4), Y => memorya289_4_Z);
    
    memorya218 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya25_3_Z, C
         => memorya162_2_Z, D => memorya474_5_Z, Y => 
        memorya218_Z);
    
    memory_memory_0_0_sr_RNO_223 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_299, B => memoryro_171, C => 
        memorya299_Z, D => memorya171_Z, Y => memoryror_85);
    
    memorya74 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya42_0_Z, B => memorya68_4_Z, C => 
        memorya41_3_Z, D => memorya84_2_Z, Y => memorya74_Z);
    
    memorya511 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya54_2_Z, B => InternalAddr2Memory(8), C
         => memorya463_5_Z, D => memorya482_2_Z, Y => 
        memorya511_Z);
    
    memorya422 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_1_Z, B => InternalAddr2Memory(6), 
        C => memorya358_6_Z, D => memorya434_2_Z, Y => 
        memorya422_Z);
    
    memorya212 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya116_1_Z, 
        C => memorya340_6_Z, D => memorya482_2_Z, Y => 
        memorya212_Z);
    
    memory_memory_0_0_sr_RNO_88 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_82, B => memoryro_274, C => 
        memorya274_Z, D => memorya82_Z, Y => memoryror_208);
    
    memoryrff_412 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_412, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_412);
    
    memoryrff_394 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_394, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_394);
    
    memorya206 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya77_2_Z, B => memorya102_1_Z, C => 
        memorya199_0_Z, D => memorya162_2_Z, Y => memorya206_Z);
    
    memory_memory_0_0_sr_RNO_383 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya20_6_Z, B => memorya116_1_Z, C => 
        memorya20_0_Z, Y => memorya20);
    
    memorya255 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya54_2_Z, B => InternalAddr2Memory(8), C
         => memorya463_5_Z, D => memorya482_2_Z, Y => 
        memorya255_Z);
    
    memoryrff_503_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya503_Z, B => WriteEnable, Y => 
        memorywre_503);
    
    memoryrff_502_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya502_Z, B => WriteEnable, Y => 
        memorywre_502);
    
    memoryrff_158 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_158, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_158);
    
    memoryrff_446 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_446, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_446);
    
    memorya245 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya54_2_Z, B => memorya117_1_Z, C => 
        memorya482_2_Z, D => memorya5_0_Z, Y => memorya245_Z);
    
    memoryrff_414 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_414, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_414);
    
    memoryrff_178 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_178, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_178);
    
    memoryrff_321_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya321_Z, B => WriteEnable, Y => 
        memorywre_321);
    
    memoryrff_257 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_257, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_257);
    
    memorya380 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya68_2_Z, C
         => memorya368_2_Z, D => memorya380_5_Z, Y => 
        memorya380_Z);
    
    memoryrff_280_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya280_Z, B => WriteEnable, Y => 
        memorywre_280);
    
    memorya478 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya370_3_Z, 
        C => memorya126_5_Z, D => memorya482_2_Z, Y => 
        memorya478_Z);
    
    memorya374 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_3_Z, B => InternalAddr2Memory(7), 
        C => memorya118_5_Z, D => memorya368_2_Z, Y => 
        memorya374_Z);
    
    memoryrff_98 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_98, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_98);
    
    memorya504_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya498_3_Z, B => memorya68_2_Z, Y => 
        memorya504_6_Z);
    
    memorya20_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(3), Y => memorya20_3_Z);
    
    memoryrff_277 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_277, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_277);
    
    memoryrff_318_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya318_Z, B => WriteEnable, Y => 
        memorywre_318);
    
    memorya344_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya25_3_Z, B => memorya68_2_Z, Y => 
        memorya344_6_Z);
    
    memorya326 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya102_1_Z, 
        C => memorya326_6_Z, D => memorya368_2_Z, Y => 
        memorya326_Z);
    
    memorya153 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya121_1_Z, B => InternalAddr2Memory(8), 
        C => memorya280_6_Z, D => memorya403_2_Z, Y => 
        memorya153_Z);
    
    memorya72 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya77_2_Z, B => memorya41_3_Z, C => 
        memorya20_0_Z, D => memorya68_4_Z, Y => memorya72_Z);
    
    memoryrff_156_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya156_Z, B => WriteEnable, Y => 
        memorywre_156);
    
    memorya2 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya2_0_Z, B => InternalAddr2Memory(8), C
         => memorya368_4_Z, D => memorya4_6_Z, Y => memorya2_Z);
    
    memoryrff_136_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya395_2_Z, B => WriteEnable, C => 
        memorya264_6_Z, D => memorya20_0_Z, Y => memorywre_136);
    
    memorya143 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya143_0_Z, B => memorya273_4_Z, C => 
        memorya463_5_Z, Y => memorya143_Z);
    
    memory_memory_0_0_sr_RNO_194 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_129, B => memoryro_257, C => 
        memorya257_Z, D => memorya129_Z, Y => memoryror_129);
    
    memoryrff_312 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_312, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_312);
    
    memory_memory_0_0_sr_RNO_151 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_356, B => memoryro_164, C => 
        memorya356_Z, D => memorya164_Z, Y => memoryror_169);
    
    memorya294 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_1_Z, B => InternalAddr2Memory(7), 
        C => memorya294_6_Z, D => memorya305_2_Z, Y => 
        memorya294_Z);
    
    memorya175 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya289_4_Z, 
        C => memorya434_2_Z, D => memorya463_5_Z, Y => 
        memorya175_Z);
    
    memoryrff_431 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_431, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_431);
    
    memorya369_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya116_2_Z, B => memorya369_1_Z, Y => 
        memorya369_5_Z);
    
    memorya168 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya45_2_Z, C
         => memorya162_2_Z, D => memorya296_6_Z, Y => 
        memorya168_Z);
    
    memorya225 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya353_1_Z, 
        C => memorya353_6_Z, D => memorya482_2_Z, Y => 
        memorya225_Z);
    
    memory_memory_0_0_sr_RNO_214 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_10, B => memoryro_394, C => 
        memorya394_Z, D => memorya10, Y => memoryror_92);
    
    memory_memory_0_0_sr_RNO_372 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya315_5_Z, B => memorya111_0_Z, C => 
        memorya211_3_Z, Y => memorya251);
    
    memoryrff_360 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_360, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_360);
    
    memoryrff_231 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_231, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_231);
    
    memoryrff_202 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_202, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_202);
    
    memoryrff_288 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_288, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_288);
    
    memoryrff_316 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_316, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_316);
    
    memory_memory_0_0_sr_RNO_164 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_185, B => memoryro_393, C => 
        memorya393_Z, D => memorya185_Z, Y => memoryror_157);
    
    memorya66 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya68_4_Z, B => memorya10_0_Z, C => 
        memorya68_3_Z, D => memorya66_1_Z, Y => memorya66_Z);
    
    memorya488 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(4), B => memorya45_2_Z, C
         => memorya376_6_Z, D => memorya482_2_Z, Y => 
        memorya488_Z);
    
    memorya384 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_2_Z, B => InternalAddr2Memory(6), C
         => memorya320_6_Z, D => memorya498_3_Z, Y => 
        memorya384_Z);
    
    memorya117_3 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(1), Y => memorya117_3_Z);
    
    memory_memory_0_0_sr_RNO_115 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_227, B => memoryro_355, C => 
        memorya355_Z, D => memorya227_Z, Y => memoryror_232);
    
    memorya63 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya52_4, B => memorya63_0, C => 
        memorya463_5_Z, Y => memorya63_Z);
    
    memorya52_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya116_1_Z, B => InternalAddr2Memory(8), 
        Y => memorya52_0_Z);
    
    memorya298_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya289_4_Z, B => memorya354_3_Z, Y => 
        memorya298_6_Z);
    
    memorya495 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya116_2_Z, B => InternalAddr2Memory(4), 
        C => memorya463_5_Z, D => memorya498_3_Z, Y => 
        memorya495_Z);
    
    memory_memory_0_0_sr_RNO_73 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_9, B => memoryror_10, C => 
        memoryror_11, D => memoryror_8, Y => memoryror_386);
    
    memory_memory_0_0_sr_RNO_315 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_162, B => memoryro_482, C => 
        memorya482_Z, D => memorya162_Z, Y => memoryror_32);
    
    memory_memory_0_0_sr_RNO_211 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_437, B => memoryro_133, C => 
        memorya437_Z, D => memorya133_Z, Y => memoryror_187);
    
    \memory_memory_0_0_OLDA_RNI8LU31[21]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(21), C => 
        memory_memory_0_0_OLDA_Z(21), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(21));
    
    memoryrff_417 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_417, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_417);
    
    memoryrff_283_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya283_Z, B => WriteEnable, Y => 
        memorywre_283);
    
    memoryrff_24_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya24_Z, B => WriteEnable, Y => 
        memorywre_24);
    
    memorya463 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya463_4_Z, B => InternalAddr2Memory(5), 
        C => memorya463_5_Z, D => memorya482_2_Z, Y => 
        memorya463_Z);
    
    memoryrff_174_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya174_Z, B => WriteEnable, Y => 
        memorywre_174);
    
    memorya369_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya369_3_Z, B => memorya368_4_Z, Y => 
        memorya369_6_Z);
    
    memorya162 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya162_2_Z, B => memorya289_6_Z, C => 
        InternalAddr2Memory(8), D => memorya354_1_Z, Y => 
        memorya162_Z);
    
    memory_memory_0_0_sr_RNO_210 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_180, B => memoryro_372, C => 
        memorya372_Z, D => memorya180_Z, Y => memoryror_185);
    
    memorya433 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya369_1_Z, B => InternalAddr2Memory(6), 
        C => memorya369_6_Z, D => memorya434_2_Z, Y => 
        memorya433_Z);
    
    memoryrff_80_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya86_2_Z, B => WriteEnable, C => 
        memorya83_6_Z, D => memorya20_0_Z, Y => memorywre_80);
    
    memorya50 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya52_2_Z, B => memorya51_6_Z, C => 
        InternalAddr2Memory(8), D => memorya370_1_Z, Y => 
        memorya50_Z);
    
    memorya185 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya193_2_Z, B => memorya121_5_Z, C => 
        InternalAddr2Memory(8), D => memorya312_4_Z, Y => 
        memorya185_Z);
    
    memorya132 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya273_4_Z, B => memorya20_0_Z, C => 
        memorya68_3_Z, D => memorya391_2_Z, Y => memorya132_Z);
    
    memoryrff_445 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_445, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_445);
    
    memoryrff_247_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya167_3_Z, C => 
        memorya503_5_Z, D => memorya111_0_Z, Y => memorywre_247);
    
    memorya105_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya102_4_Z, B => memorya57_3_Z, Y => 
        memorya105_6_Z);
    
    memoryrff_190 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_190, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_190);
    
    memoryrff_500_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya500_Z, B => WriteEnable, Y => 
        memorywre_500);
    
    memoryrff_171_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya171_Z, B => WriteEnable, Y => 
        memorywre_171);
    
    memoryrff_100_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya100_Z, B => WriteEnable, Y => 
        memorywre_100);
    
    memoryrff_451_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya451_Z, B => WriteEnable, Y => 
        memorywre_451);
    
    memorya279 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya487_4_Z, 
        C => memorya273_4_Z, D => memorya503_5_Z, Y => 
        memorya279_Z);
    
    memoryrff_431_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya431_Z, B => WriteEnable, Y => 
        memorywre_431);
    
    memoryrff_112 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_112, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_112);
    
    memoryrff_98_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya98_Z, B => WriteEnable, Y => 
        memorywre_98);
    
    memoryrff_38_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya38_Z, B => WriteEnable, Y => 
        memorywre_38);
    
    memoryrff_275_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya275_Z, B => WriteEnable, Y => 
        memorywre_275);
    
    memorya51_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya52_4, B => memorya368_4_Z, Y => 
        memorya51_6_Z);
    
    memorya267 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya264_1_Z, B => memorya264_6_Z, C => 
        InternalAddr2Memory(7), D => memorya379_1_Z, Y => 
        memorya267_Z);
    
    memoryrff_90 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_90, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_90);
    
    memoryrff_54_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya54_Z, B => WriteEnable, Y => 
        memorywre_54);
    
    memoryrff_175_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya175_Z, B => WriteEnable, Y => 
        memorywre_175);
    
    memorya237 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya45_2_Z, B => memorya117_1_Z, C => 
        memorya482_2_Z, D => memorya236_0_Z, Y => memorya237_Z);
    
    memoryrff_354 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_354, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_354);
    
    memorya345_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya86_2_Z, B => memorya121_1_Z, Y => 
        memorya345_5_Z);
    
    memory_memory_0_0_sr_RNO_380 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya84_2_Z, B => memorya124_0_Z, C => 
        memorya380_5_Z, Y => memorya124);
    
    memorya280_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya273_4_Z, B => memorya57_3_Z, Y => 
        memorya280_6_Z);
    
    memorya256 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_3_Z, B => InternalAddr2Memory(7), C
         => memorya376_6_Z, D => memorya273_4_Z, Y => 
        memorya256_Z);
    
    memory_memory_0_0_sr_RNO_352 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya315_5_Z, B => memorya111_0_Z, C => 
        memorya121_4_Z, Y => memorya123);
    
    memoryrff_264_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya264_Z, B => WriteEnable, Y => 
        memorywre_264);
    
    memoryrff_272_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya272_Z, B => WriteEnable, Y => 
        memorywre_272);
    
    memoryrff_143_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya143_Z, B => WriteEnable, Y => 
        memorywre_143);
    
    memoryrff_97_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya97_Z, B => WriteEnable, Y => 
        memorywre_97);
    
    memoryrff_37_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya37_Z, B => WriteEnable, Y => 
        memorywre_37);
    
    memoryrff_374 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_374, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_374);
    
    memorya246 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya102_3_Z, 
        C => memorya118_5_Z, D => memorya482_2_Z, Y => 
        memorya246_Z);
    
    memory_memory_0_0_sr_RNO_236 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_73, B => memoryro_329, C => 
        memorya329_Z, D => memorya73_Z, Y => memoryror_77);
    
    memoryrff_409_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya409_Z, B => WriteEnable, Y => 
        memorywre_409);
    
    memorya476 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya86_2_Z, B => memorya504_6_Z, C => 
        InternalAddr2Memory(5), D => memorya364_1_Z, Y => 
        memorya476_Z);
    
    memorya367 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya463_4_Z, 
        C => memorya116_2_Z, D => memorya463_5_Z, Y => 
        memorya367_Z);
    
    memoryrff_345_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya345_Z, B => WriteEnable, Y => 
        memorywre_345);
    
    memorya337 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya368_2_Z, B => memorya336_6_Z, C => 
        InternalAddr2Memory(7), D => memorya369_1_Z, Y => 
        memorya337_Z);
    
    memorya289_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya289_4_Z, B => memorya368_4_Z, Y => 
        memorya289_6_Z);
    
    memory_memory_0_0_sr_RNO_42 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_155, B => memoryror_153, C => 
        memoryror_152, D => memoryror_154, Y => memoryror_422);
    
    memoryrff_21 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_21, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_21);
    
    memoryrff_187 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_187, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_187);
    
    memoryrff_214 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_214, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_214);
    
    memorya86_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya86_2_Z, B => memorya102_1_Z, Y => 
        memorya86_5_Z);
    
    memoryrff_208 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_208, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_208);
    
    memoryrff_148 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_148, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_148);
    
    memory_memory_0_0_sr_RNO_117 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_414, B => memoryro_78, C => 
        memorya414_Z, D => memorya78_Z, Y => memoryror_199);
    
    memorya289 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya353_1_Z, B => InternalAddr2Memory(7), 
        C => memorya289_6_Z, D => memorya369_3_Z, Y => 
        memorya289_Z);
    
    memoryrff_297_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya297_Z, B => WriteEnable, Y => 
        memorywre_297);
    
    memoryrff_383 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_383, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_383);
    
    memoryrff_224_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya224_Z, B => WriteEnable, Y => 
        memorywre_224);
    
    memorya52_2 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(0), Y => memorya52_2_Z);
    
    memoryrff_330 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_330, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_330);
    
    memoryrff_247 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_247, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_247);
    
    memorya226 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya354_1_Z, 
        C => memorya354_6_Z, D => memorya482_2_Z, Y => 
        memorya226_Z);
    
    memoryrff_421 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_421, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_421);
    
    memory_memory_0_0_sr_RNO_279 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_295, B => memoryro_39, C => 
        memorya295_Z, D => memorya39_Z, Y => memoryror_62);
    
    memory_memory_0_0_sr_RNO_275 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_387, B => memoryro_115, C => 
        memorya387_Z, D => memorya115_Z, Y => memoryror_120);
    
    \memory_memory_0_0_OLDA[19]\ : SLE
      port map(D => \InternalDataFromMem\(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(19));
    
    memoryrff_109_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya109_Z, B => WriteEnable, Y => 
        memorywre_109);
    
    memoryrff_221 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_221, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_221);
    
    memorya12_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya364_1_Z, B => InternalAddr2Memory(8), 
        Y => memorya12_0_Z);
    
    memorya102_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya116_2_Z, B => memorya102_1_Z, Y => 
        memorya102_5_Z);
    
    memorya486 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_3_Z, B => InternalAddr2Memory(4), 
        C => memorya102_5_Z, D => memorya498_3_Z, Y => 
        memorya486_Z);
    
    memory_memory_0_0_sr_RNO_29 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_206, B => memoryror_205, C => 
        memoryror_207, D => memoryror_204, Y => memoryror_435);
    
    memorya31 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya31_0_Z, C
         => memorya463_5_Z, D => memorya52_4, Y => memorya31_Z);
    
    memorya391_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(2), Y => memorya391_2_Z);
    
    memoryrff_510 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_510, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_510);
    
    memoryrff_357_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya357_Z, B => WriteEnable, Y => 
        memorywre_357);
    
    memoryrff_337_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya337_Z, B => WriteEnable, Y => 
        memorywre_337);
    
    memoryrff_193_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya193_Z, B => WriteEnable, Y => 
        memorywre_193);
    
    memorya68_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(2), Y => memorya68_1_Z);
    
    memoryrff_26_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya26_Z, B => WriteEnable, Y => 
        memorywre_26);
    
    memoryrff_395_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya395_Z, B => WriteEnable, Y => 
        memorywre_395);
    
    memoryrff_464_RNO : CFG3
      generic map(INIT => x"80")

      port map(A => memorya464_0_Z, B => WriteEnable, C => 
        memorya368_6_Z, Y => memorywre_464);
    
    memory_memory_0_0_sr_RNO_70 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_53, B => memoryror_55, C => 
        memoryror_54, D => memoryror_52, Y => memoryror_397);
    
    \memory_memory_0_0_OLDA_RNICOT31[16]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(16), C => 
        memory_memory_0_0_OLDA_Z(16), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(16));
    
    memory_memory_0_0_en : SLE
      port map(D => dout_1_sqmuxa_Z, CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => memory_memory_0_0_en_Z);
    
    memorya353_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya57_3_Z, B => memorya68_3_Z, Y => 
        memorya353_6_Z);
    
    memorya128_0 : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory(8), B => memorya57_3_Z, C
         => memorya162_2_Z, Y => memorya128_0_Z);
    
    memory_memory_0_0_sr_RNO_26 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_238, B => memoryror_236, C => 
        memoryror_237, D => memoryror_239, Y => memoryror_443);
    
    memorya55 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya55_0_Z, C
         => memorya503_5_Z, D => memorya52_4, Y => memorya55_Z);
    
    memorya46 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya46_3_Z, C
         => memorya52_4, D => memorya110_5_Z, Y => memorya46_Z);
    
    memory_memory_0_0_sr_RNO_329 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_285, B => memoryro_45, C => 
        memorya285_Z, D => memorya45_Z, Y => memoryror_22);
    
    memorya43 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya41_3_Z, C
         => memorya52_4, D => memorya299_5_Z, Y => memorya43_Z);
    
    memorya361 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya121_1_Z, 
        C => memorya116_2_Z, D => memorya361_6_Z, Y => 
        memorya361_Z);
    
    memorya54 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya102_3_Z, 
        C => memorya52_4, D => memorya118_5_Z, Y => memorya54_Z);
    
    memorya30_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(0), Y => memorya30_3_Z);
    
    memorya331 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya4_3_Z, B => InternalAddr2Memory(7), C
         => memorya331_5_Z, D => memorya379_4_Z, Y => 
        memorya331_Z);
    
    memorya121_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(0), Y => memorya121_1_Z);
    
    memoryrff_150 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_150, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_150);
    
    memory_memory_0_0_sr_RNO_63 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_103, B => memoryror_102, C => 
        memoryror_100, D => memoryror_101, Y => memoryror_409);
    
    memoryrff_41 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_41, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_41);
    
    memorya191 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(7), C => memorya63_0, D => 
        memorya463_5_Z, Y => memorya191_Z);
    
    memoryrff_170 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_170, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_170);
    
    memorya85 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya84_3_Z, C
         => memorya68_4_Z, D => memorya213_5_Z, Y => memorya85_Z);
    
    memory_memory_0_0_sr_RNO_146 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_213, B => memoryro_485, C => 
        memorya485_Z, D => memorya213_Z, Y => memoryror_251);
    
    memoryrff_510_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya510_Z, B => WriteEnable, Y => 
        memorywre_510);
    
    memorya326_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya4_3_Z, B => memorya102_3_Z, Y => 
        memorya326_6_Z);
    
    memoryrff_424_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya424_Z, B => WriteEnable, Y => 
        memorywre_424);
    
    memoryrff_215 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_215, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_215);
    
    memorya84 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya84_2_Z, B => memorya84_3_Z, C => 
        memorya68_4_Z, D => memorya52_0_Z, Y => memorya84_Z);
    
    memory_memory_0_0_sr_RNO_324 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_31, B => memoryro_287, C => 
        memorya287_Z, D => memorya31_Z, Y => memoryror_19);
    
    memoryrff_110_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya110_Z, B => WriteEnable, Y => 
        memorywre_110);
    
    memoryrff_107 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_107, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_107);
    
    \memory_memory_0_0_OLDA[17]\ : SLE
      port map(D => \InternalDataFromMem\(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(17));
    
    memoryrff_457_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya457_Z, B => WriteEnable, Y => 
        memorywre_457);
    
    memorya261 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya273_4_Z, B => memorya68_3_Z, C => 
        memorya261_0_Z, D => memorya369_3_Z, Y => memorya261_Z);
    
    memorya257_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya273_4_Z, B => memorya68_3_Z, Y => 
        memorya257_6_Z);
    
    memoryrff_56_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya56_Z, B => WriteEnable, Y => 
        memorywre_56);
    
    memoryrff_437_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya437_Z, B => WriteEnable, Y => 
        memorywre_437);
    
    memorya231 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya482_2_Z, B => memorya227_0_Z, C => 
        memorya487_5_Z, Y => memorya231_Z);
    
    memory_memory_0_0_sr_RNO_259 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_283, B => memoryro_155, C => 
        memorya283_Z, D => memorya155_Z, Y => memoryror_101);
    
    memory_memory_0_0_sr_RNO_255 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_401, B => memoryro_33, C => 
        memorya401_Z, D => memorya33_Z, Y => memoryror_97);
    
    memorya107 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya67_2_Z, C
         => memorya102_4_Z, D => memorya299_5_Z, Y => 
        memorya107_Z);
    
    memoryrff_16 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_16, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_16);
    
    memorya412 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya29_3_Z, B => InternalAddr2Memory(6), C
         => memorya156_5_Z, D => memorya370_3_Z, Y => 
        memorya412_Z);
    
    memory_memory_0_0_sr_RNO_326 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_81, B => memoryro_497, C => 
        memorya497, D => memorya81_Z, Y => memoryror_17);
    
    memorya52 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya52_2_Z, B => memorya84_3_Z, C => 
        memorya52_4, D => memorya52_0_Z, Y => memorya52_Z);
    
    memorya390 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya102_1_Z, 
        C => memorya326_6_Z, D => memorya498_3_Z, Y => 
        memorya390_Z);
    
    memoryrff_303 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_303, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_303);
    
    memoryrff_381 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_381, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_381);
    
    memory_memory_0_0_sr_RNO_111 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_360, B => memoryro_152, C => 
        memorya360_Z, D => memorya152_Z, Y => memoryror_239);
    
    memoryrff_501_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya501_Z, B => WriteEnable, Y => 
        memorywre_501);
    
    memoryrff_419_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya419_Z, B => WriteEnable, Y => 
        memorywre_419);
    
    memoryrff_40_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya40_Z, B => WriteEnable, Y => 
        memorywre_40);
    
    memory_memory_0_0_sr_RNO_206 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_0, B => memoryro_304, C => 
        memorya304_Z, D => memorya0, Y => memoryror_178);
    
    memoryrff_63_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya63_Z, B => WriteEnable, Y => 
        memorywre_63);
    
    memoryrff_276_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya276_Z, B => WriteEnable, Y => 
        memorywre_276);
    
    memoryrff_365 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_365, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_365);
    
    memoryrff_344 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_344, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_344);
    
    memorya508 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(1), B => memorya370_3_Z, 
        C => memorya380_5_Z, D => memorya482_2_Z, Y => 
        memorya508_Z);
    
    memoryrff_185 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_185, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_185);
    
    memorya82 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya84_2_Z, B => memorya83_6_Z, C => 
        InternalAddr2Memory(8), D => memorya370_1_Z, Y => 
        memorya82_Z);
    
    \memory_memory_0_0_OLDA_RNIBNT31[15]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(15), C => 
        memory_memory_0_0_OLDA_Z(15), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(15));
    
    memorya41_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(2), Y => memorya41_3_Z);
    
    memorya316 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya316_4_Z, 
        C => memorya370_3_Z, D => memorya380_5_Z, Y => 
        memorya316_Z);
    
    \memory_memory_0_0_OLDA[11]\ : SLE
      port map(D => \InternalDataFromMem\(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(11));
    
    memoryrff_358_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya358_Z, B => WriteEnable, Y => 
        memorywre_358);
    
    memory_memory_0_0_sr_RNO_148 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_291, B => memoryro_163, C => 
        memorya291_Z, D => memorya163_Z, Y => memoryror_168);
    
    memoryrff_338_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya338_Z, B => WriteEnable, Y => 
        memorywre_338);
    
    memorya71 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_3_Z, B => InternalAddr2Memory(8), C
         => memorya455_5_Z, D => memorya68_4_Z, Y => memorya71_Z);
    
    memoryrff_344_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya344_Z, B => WriteEnable, Y => 
        memorywre_344);
    
    memoryrff_369 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_369, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_369);
    
    memorya294_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya289_4_Z, B => memorya102_3_Z, Y => 
        memorya294_6_Z);
    
    memorya25_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(2), Y => memorya25_3_Z);
    
    memory_memory_0_0_sr_RNO_93 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_245, B => memoryro_453, C => 
        memorya453_Z, D => memorya245_Z, Y => memoryror_219);
    
    memoryrff_320 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_320, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_320);
    
    memorya360_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya68_2_Z, B => memorya41_3_Z, Y => 
        memorya360_6_Z);
    
    memoryrff_5 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_5, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_5);
    
    memoryrff_25_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya25_Z, B => WriteEnable, Y => 
        memorywre_25);
    
    memorya302 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya289_4_Z, B => InternalAddr2Memory(7), 
        C => memorya110_5_Z, D => memorya370_3_Z, Y => 
        memorya302_Z);
    
    memorya193_2 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(1), Y => memorya193_2_Z);
    
    memoryrff_86 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_86, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_86);
    
    memoryrff_491 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_491, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_491);
    
    memorya215 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya211_0_Z, B => memorya482_2_Z, C => 
        memorya503_5_Z, Y => memorya215_Z);
    
    \memory_memory_0_0_OLDA_RNINOUT[2]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(2), C => 
        memory_memory_0_0_OLDA_Z(2), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(2));
    
    memorya109 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya117_1_Z, B => memorya45_2_Z, C => 
        memorya102_4_Z, D => memorya93_0, Y => memorya109_Z);
    
    memorya154_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya403_2_Z, B => memorya362_1_Z, Y => 
        memorya154_5_Z);
    
    memory_memory_0_0_sr_RNO_184 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_395, B => memoryro_123, C => 
        memorya395_Z, D => memorya123, Y => memoryror_133);
    
    memoryrff_119_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya116_4_Z, C => 
        memorya503_5_Z, D => memorya111_0_Z, Y => memorywre_119);
    
    memorya498 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(3), B => memorya370_1_Z, 
        C => memorya116_2_Z, D => memorya498_6_Z, Y => 
        memorya498_Z);
    
    memorya394 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya362_1_Z, 
        C => memorya202_6_Z, D => memorya498_3_Z, Y => 
        memorya394_Z);
    
    memoryrff_506 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_506, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_506);
    
    memoryrff_291 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_291, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_291);
    
    memoryrff_164_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya164_Z, B => WriteEnable, Y => 
        memorywre_164);
    
    memorya467 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya379_1_Z, 
        C => memorya86_2_Z, D => memorya435_6_Z, Y => 
        memorya467_Z);
    
    memorya437 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya84_3_Z, C
         => memorya373_5_Z, D => memorya498_3_Z, Y => 
        memorya437_Z);
    
    memory_memory_0_0_sr_RNO_33 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_255, B => memoryror_252, C => 
        memoryror_254, D => memoryror_253, Y => memoryror_447);
    
    memory_memory_0_0_sr_RNO_173 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_340, B => memoryro_148, C => 
        memorya340_Z, D => memorya148_Z, Y => memoryror_153);
    
    memory_memory_0_0_sr_RNO_132 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_241, B => memoryro_369, C => 
        memorya369_Z, D => memorya241, Y => memoryror_241);
    
    memorya502 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(3), B => memorya370_3_Z, 
        C => memorya118_5_Z, D => memorya482_2_Z, Y => 
        memorya502_Z);
    
    memorya409 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya121_1_Z, B => InternalAddr2Memory(6), 
        C => memorya345_6_Z, D => memorya403_2_Z, Y => 
        memorya409_Z);
    
    memorya303 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya289_4_Z, 
        C => memorya305_2_Z, D => memorya463_5_Z, Y => 
        memorya303_Z);
    
    memorya166 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_1_Z, B => InternalAddr2Memory(8), 
        C => memorya294_6_Z, D => memorya434_2_Z, Y => 
        memorya166_Z);
    
    memorya113 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya57_3_Z, C
         => memorya116_4_Z, D => memorya369_5_Z, Y => 
        memorya113_Z);
    
    memoryrff_507_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya507_Z, B => WriteEnable, Y => 
        memorywre_507);
    
    memoryrff_161_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya161_Z, B => WriteEnable, Y => 
        memorywre_161);
    
    memorya68_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(3), Y => memorya68_3_Z);
    
    memorya276_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya116_1_Z, B => InternalAddr2Memory(7), 
        Y => memorya276_0_Z);
    
    memorya195 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_1_Z, B => InternalAddr2Memory(8), 
        C => memorya320_6_Z, D => memorya482_2_Z, Y => 
        memorya195_Z);
    
    memorya193_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(0), Y => memorya193_1_Z);
    
    memoryrff_55_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya55_Z, B => WriteEnable, Y => 
        memorywre_55);
    
    memoryrff_483 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_483, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_483);
    
    memoryrff_480 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_480, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_480);
    
    memoryrff_265_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya265_Z, B => WriteEnable, Y => 
        memorywre_265);
    
    memorya160 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya368_4_Z, B => memorya289_4_Z, C => 
        memorya434_2_Z, D => memorya20_0_Z, Y => memorya160_Z);
    
    memoryrff_165_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya165_Z, B => WriteEnable, Y => 
        memorywre_165);
    
    memoryrff_124_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya124_0_Z, B => memorya380_5_Z, C => 
        WriteEnable, D => memorya84_2_Z, Y => memorywre_124);
    
    memorya130 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya273_4_Z, B => memorya10_0_Z, C => 
        memorya68_3_Z, D => memorya386_1_Z, Y => memorya130_Z);
    
    memorya379_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(1), Y => memorya379_1_Z);
    
    memorya354_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(2), Y => memorya354_3_Z);
    
    memoryrff_68 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_68, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_68);
    
    memoryrff_394_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya394_Z, B => WriteEnable, Y => 
        memorywre_394);
    
    memoryrff_262_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya262_Z, B => WriteEnable, Y => 
        memorywre_262);
    
    memory_memory_0_0_sr_RNO_312 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_47, B => memoryro_303, C => 
        memorya303_Z, D => memorya47_Z, Y => memoryror_35);
    
    memoryrff_509 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_509, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_509);
    
    memory_memory_0_0_sr_RNO_60 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_111, B => memoryror_110, C => 
        memoryror_108, D => memoryror_109, Y => memoryror_411);
    
    memoryrff_503 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_503, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_503);
    
    memoryrff_301 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_301, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_301);
    
    memory_memory_0_0_sr_RNO_14 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_411, B => memoryror_410, C => 
        memoryror_408, D => memoryror_409, Y => memoryror_486);
    
    memoryrff_184 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_184, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_184);
    
    memoryrff_121_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya121_Z, B => WriteEnable, Y => 
        memorywre_121);
    
    \memory_memory_0_0_OLDA[9]\ : SLE
      port map(D => \InternalDataFromMem\(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(9));
    
    memoryrff_318 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_318, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_318);
    
    memoryrff_13 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_13, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_13);
    
    memoryrff_176_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya176_Z, B => WriteEnable, Y => 
        memorywre_176);
    
    memoryrff_140 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_140, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_140);
    
    memoryrff_105 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_105, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_105);
    
    memorya157 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya273_4_Z, 
        C => memorya193_2_Z, D => memorya381_5_Z, Y => 
        memorya157_Z);
    
    memoryrff_225_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya225_Z, B => WriteEnable, Y => 
        memorywre_225);
    
    memoryrff_125_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya125_Z, B => WriteEnable, Y => 
        memorywre_125);
    
    memorya147 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_1_Z, B => InternalAddr2Memory(8), 
        C => memorya273_6_Z, D => memorya403_2_Z, Y => 
        memorya147_Z);
    
    memoryrff_38 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_38, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_38);
    
    memoryrff_335 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_335, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_335);
    
    memorya503 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya116_2_Z, B => InternalAddr2Memory(3), 
        C => memorya503_5_Z, D => memorya498_3_Z, Y => 
        memorya503_Z);
    
    memoryrff_222_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya222_Z, B => WriteEnable, Y => 
        memorywre_222);
    
    memory_memory_0_0_sr_RNO_153 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_239, B => memoryro_431, C => 
        memorya431_Z, D => memorya239_Z, Y => memoryror_163);
    
    memoryrff_405_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya405_Z, B => WriteEnable, Y => 
        memorywre_405);
    
    memoryrff_511_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya511_Z, B => WriteEnable, Y => 
        memorywre_511);
    
    memorya299 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya289_4_Z, B => InternalAddr2Memory(7), 
        C => memorya299_5_Z, D => memorya379_4_Z, Y => 
        memorya299_Z);
    
    memoryrff_339 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_339, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_339);
    
    memoryrff_147_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya147_Z, B => WriteEnable, Y => 
        memorywre_147);
    
    memory_memory_0_0_sr_RNO_277 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_313, B => memoryro_57, C => 
        memorya313_Z, D => memorya57_Z, Y => memoryror_61);
    
    memory_memory_0_0_sr_RNO_238 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_26, B => memoryro_410, C => 
        memorya410_Z, D => memorya26_Z, Y => memoryror_76);
    
    memoryrff_64_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya64_Z, B => WriteEnable, Y => 
        memorywre_64);
    
    memoryrff_418 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_418, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_418);
    
    \memory_memory_0_0_OLDA[28]\ : SLE
      port map(D => \InternalDataFromMem\(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(28));
    
    memoryrff_83 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_83, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_83);
    
    memoryrff_508 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_508, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_508);
    
    memorya127 : CFG4
      generic map(INIT => x"2000")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(7), C => memorya63_0, D => 
        memorya463_5_Z, Y => memorya127_Z);
    
    memorya500 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(3), B => memorya116_1_Z, 
        C => memorya116_2_Z, D => memorya504_6_Z, Y => 
        memorya500_Z);
    
    memory_memory_0_0_sr_RNO_1 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_490, B => memoryror_489, C => 
        memoryror_488, D => memoryror_491, Y => memoryror_506);
    
    memoryrff_451 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_451, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_451);
    
    memoryrff_390 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_390, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_390);
    
    memorya352 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya116_2_Z, 
        C => memorya353_6_Z, D => memorya370_3_Z, Y => 
        memorya352_Z);
    
    memorya216 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya125_2_Z, 
        C => memorya344_6_Z, D => memorya482_2_Z, Y => 
        memorya216_Z);
    
    memorya496 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(3), B => memorya54_2_Z, C
         => memorya376_6_Z, D => memorya482_2_Z, Y => 
        memorya496_Z);
    
    memoryrff_482_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya482_Z, B => WriteEnable, Y => 
        memorywre_482);
    
    memoryrff_249_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya249_Z, B => WriteEnable, Y => 
        memorywre_249);
    
    memorya159 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya273_4_Z, 
        C => memorya403_2_Z, D => memorya463_5_Z, Y => 
        memorya159_Z);
    
    memory_memory_0_0_sr_RNO_90 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_336, B => memoryro_96, C => 
        memorya336_Z, D => memorya96_Z, Y => memoryror_210);
    
    memorya376_6 : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(8), C => memorya57_3_Z, Y => 
        memorya376_6_Z);
    
    memorya342 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya86_2_Z, B => memorya342_6_Z, C => 
        InternalAddr2Memory(7), D => memorya102_1_Z, Y => 
        memorya342_Z);
    
    memoryrff_471 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_471, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_471);
    
    memoryrff_286 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_286, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_286);
    
    memoryrff_251 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_251, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_251);
    
    memorya149 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya84_3_Z, B => InternalAddr2Memory(8), C
         => memorya149_5_Z, D => memorya273_4_Z, Y => 
        memorya149_Z);
    
    memoryrff_403 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_403, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_403);
    
    memoryrff_400 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_400, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_400);
    
    memoryrff_271 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_271, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_271);
    
    \memory_memory_0_0_OLDA_RNIUVUT[9]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(9), C => 
        memory_memory_0_0_OLDA_Z(9), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(9));
    
    memorya459 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya41_3_Z, B => InternalAddr2Memory(5), C
         => memorya331_5_Z, D => memorya498_3_Z, Y => 
        memorya459_Z);
    
    memorya353 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya353_1_Z, B => InternalAddr2Memory(7), 
        C => memorya353_6_Z, D => memorya368_2_Z, Y => 
        memorya353_Z);
    
    memoryrff_471_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya471_Z, B => WriteEnable, Y => 
        memorywre_471);
    
    memorya449 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya193_1_Z, 
        C => memorya353_6_Z, D => memorya498_3_Z, Y => 
        memorya449_Z);
    
    memorya343 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya20_3_Z, C
         => memorya368_2_Z, D => memorya503_5_Z, Y => 
        memorya343_Z);
    
    memoryrff_60 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_60, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_60);
    
    memory_memory_0_0_sr_RNO_30 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_195, B => memoryror_192, C => 
        memoryror_194, D => memoryror_193, Y => memoryror_432);
    
    memory_memory_0_0_sr_RNO_102 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_353, B => memoryro_225, C => 
        memorya353_Z, D => memorya225_Z, Y => memoryror_225);
    
    memorya167_3 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(3), Y => memorya167_3_Z);
    
    memory_memory_0_0_sr_RNO_28 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_198, B => memoryror_199, C => 
        memoryror_196, D => memoryror_197, Y => memoryror_433);
    
    memory_memory_0_0_sr_RNO_149 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_149, B => memoryro_421, C => 
        memorya421_Z, D => memorya149_Z, Y => memoryror_171);
    
    memory_memory_0_0_sr_RNO_140 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_43, B => memoryro_491, C => 
        memorya491_Z, D => memorya43_Z, Y => memoryror_245);
    
    memoryrff_21_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya117_1_Z, C => 
        memorya21_0_Z, D => memorya20_6_Z, Y => memorywre_21);
    
    memoryrff_104 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_104, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_104);
    
    memorya322 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya66_1_Z, B => InternalAddr2Memory(7), C
         => memorya320_6_Z, D => memorya370_3_Z, Y => 
        memorya322_Z);
    
    memorya20_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya52_4, B => memorya20_3_Z, Y => 
        memorya20_6_Z);
    
    memory_memory_0_0_sr_RNO_337 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_467, B => memoryro_19, C => 
        memorya467_Z, D => memorya19_Z, Y => memoryror_24);
    
    memoryrff_197_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya197_Z, B => WriteEnable, Y => 
        memorywre_197);
    
    memorya129 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya57_3_Z, B => InternalAddr2Memory(8), C
         => memorya257_6_Z, D => memorya385_1_Z, Y => 
        memorya129_Z);
    
    memorya441_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya498_3_Z, B => memorya57_3_Z, Y => 
        memorya441_6_Z);
    
    memory_memory_0_0_sr_RNO_219 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_86, B => memoryro_342, C => 
        memorya342_Z, D => memorya86_Z, Y => memoryror_90);
    
    memory_memory_0_0_sr_RNO_215 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_89, B => memoryro_345, C => 
        memorya345_Z, D => memorya89_Z, Y => memoryror_93);
    
    memory_memory_0_0_sr_RNO_257 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_365, B => memoryro_109, C => 
        memorya365_Z, D => memorya109_Z, Y => memoryror_102);
    
    memory_memory_0_0_sr_RNO_233 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_419, B => memoryro_67, C => 
        memorya419_Z, D => memorya67_Z, Y => memoryror_72);
    
    \memory_memory_0_0_OLDA_RNI9MU31[22]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(22), C => 
        memory_memory_0_0_OLDA_Z(22), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(22));
    
    memoryrff_30 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_30, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_30);
    
    memorya429 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya45_3_Z, C
         => memorya45_5_Z, D => memorya498_3_Z, Y => memorya429_Z);
    
    memorya323 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya368_2_Z, B => memorya320_6_Z, C => 
        InternalAddr2Memory(7), D => memorya379_1_Z, Y => 
        memorya323_Z);
    
    memoryrff_260 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_260, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_260);
    
    memoryrff_299_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya299_Z, B => WriteEnable, Y => 
        memorywre_299);
    
    memoryrff_12 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_12, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_12);
    
    memorya36_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(2), Y => memorya36_1_Z);
    
    memorya482_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(6), Y => memorya482_2_Z);
    
    \memory_memory_0_0_OLDA_RNI8KT31[12]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(12), C => 
        memory_memory_0_0_OLDA_Z(12), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(12));
    
    memoryrff_266_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya266_Z, B => WriteEnable, Y => 
        memorywre_266);
    
    memoryrff_150_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya150_Z, B => WriteEnable, Y => 
        memorywre_150);
    
    memoryrff_130_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya130_Z, B => WriteEnable, Y => 
        memorywre_130);
    
    memoryrff_240_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya240_Z, B => WriteEnable, Y => 
        memorywre_240);
    
    memorya305 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya305_2_Z, B => memorya304_6_Z, C => 
        InternalAddr2Memory(7), D => memorya369_1_Z, Y => 
        memorya305_Z);
    
    memoryrff_51_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya51_Z, B => WriteEnable, Y => 
        memorywre_51);
    
    memory_memory_0_0_sr_RNO_79 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_43, B => memoryror_41, C => 
        memoryror_40, D => memoryror_42, Y => memoryror_394);
    
    memoryrff_181 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_181, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_181);
    
    memorya51 : CFG3
      generic map(INIT => x"20")

      port map(A => memorya51_6_Z, B => InternalAddr2Memory(8), C
         => memorya499_5_Z, Y => memorya51_Z);
    
    memoryrff_325 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_325, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_325);
    
    memory_memory_0_0_sr_RNO_341 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya227_0_Z, B => memorya102_5_Z, C => 
        memorya162_2_Z, Y => memorya230);
    
    memoryrff_462 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_462, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_462);
    
    memoryrff_459_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya459_Z, B => WriteEnable, Y => 
        memorywre_459);
    
    memoryrff_415_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya415_Z, B => WriteEnable, Y => 
        memorywre_415);
    
    memoryrff_439_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya439_Z, B => WriteEnable, Y => 
        memorywre_439);
    
    memoryrff_377_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya377_Z, B => WriteEnable, Y => 
        memorywre_377);
    
    memorya164 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya36_1_Z, C
         => memorya162_2_Z, D => memorya292_6_Z, Y => 
        memorya164_Z);
    
    \memory_memory_0_0_OLDA[31]\ : SLE
      port map(D => \InternalDataFromMem\(31), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(31));
    
    memoryrff_206 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_206, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_206);
    
    memoryrff_329 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_329, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_329);
    
    memoryrff_226_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya226_Z, B => WriteEnable, Y => 
        memorywre_226);
    
    memorya81 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya117_3_Z, B => memorya83_6_Z, C => 
        InternalAddr2Memory(8), D => memorya369_1_Z, Y => 
        memorya81_Z);
    
    memorya7 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya7_0_Z, B => InternalAddr2Memory(8), C
         => memorya379_1_Z, D => memorya4_6_Z, Y => memorya7_Z);
    
    memorya134 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya102_1_Z, 
        C => memorya162_2_Z, D => memorya257_6_Z, Y => 
        memorya134_Z);
    
    memory_memory_0_0_sr_RNO_76 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_39, B => memoryror_38, C => 
        memoryror_37, D => memoryror_36, Y => memoryror_393);
    
    memoryrff_66_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya66_Z, B => WriteEnable, Y => 
        memorywre_66);
    
    memoryrff_486 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_486, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_486);
    
    memoryrff_464 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_464, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_464);
    
    memoryrff_386_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya386_Z, B => WriteEnable, Y => 
        memorywre_386);
    
    memoryrff_82 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_82, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_82);
    
    memory_memory_0_0_sr_RNO_208 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_182, B => memoryro_454, C => 
        memorya454_Z, D => memorya182_Z, Y => memoryror_186);
    
    memory_memory_0_0_sr_RNO_126 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_112, B => memoryro_320, C => 
        memorya320_Z, D => memorya112_Z, Y => memoryror_194);
    
    memoryrff_350 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_350, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_350);
    
    memory_memory_0_0_sr_RNO_57 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_74, B => memoryror_72, C => 
        memoryror_75, D => memoryror_73, Y => memoryror_402);
    
    memoryrff_370 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_370, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_370);
    
    memoryrff_89_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya89_Z, B => WriteEnable, Y => 
        memorywre_89);
    
    memoryrff_362 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_362, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_362);
    
    memoryrff_243_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya243_Z, B => WriteEnable, Y => 
        memorywre_243);
    
    memorya340_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya20_3_Z, B => memorya68_2_Z, Y => 
        memorya340_6_Z);
    
    dout_1_sqmuxa : CFG2
      generic map(INIT => x"2")

      port map(A => resetn, B => WriteEnable, Y => 
        dout_1_sqmuxa_Z);
    
    memoryrff_159_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya159_Z, B => WriteEnable, Y => 
        memorywre_159);
    
    memoryrff_139_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya139_Z, B => WriteEnable, Y => 
        memorywre_139);
    
    memoryrff_290_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya290_Z, B => WriteEnable, Y => 
        memorywre_290);
    
    memory_memory_0_0_sr_RNO_296 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_404, B => memoryro_4, C => 
        memorya404_Z, D => memorya4_Z, Y => memoryror_9);
    
    memoryrff_441 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_441, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_441);
    
    memoryrff_219 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_219, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_219);
    
    memoryrff_477_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya477_Z, B => WriteEnable, Y => 
        memorywre_477);
    
    memorya434 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya370_1_Z, B => InternalAddr2Memory(6), 
        C => memorya370_6_Z, D => memorya434_2_Z, Y => 
        memorya434_Z);
    
    memory_memory_0_0_sr_RNO_87 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_344, B => memoryro_168, C => 
        memorya344_Z, D => memorya168_Z, Y => memoryror_223);
    
    memoryrff_241 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_241, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_241);
    
    memorya200 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya77_2_Z, C
         => memorya162_2_Z, D => memorya393_6_Z, Y => 
        memorya200_Z);
    
    memory_memory_0_0_sr_RNO_373 : CFG3
      generic map(INIT => x"20")

      port map(A => memorya4_6_Z, B => InternalAddr2Memory(8), C
         => memorya463_5_Z, Y => memorya15);
    
    memoryrff_508_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya508_Z, B => WriteEnable, Y => 
        memorywre_508);
    
    memoryrff_366 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_366, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_366);
    
    memoryrff_207_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya207_Z, B => WriteEnable, Y => 
        memorywre_207);
    
    memorya470 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya102_3_Z, 
        C => memorya86_5_Z, D => memorya498_3_Z, Y => 
        memorya470_Z);
    
    memory_memory_0_0_sr_RNO_128 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_198, B => memoryro_406, C => 
        memorya406_Z, D => memorya198_Z, Y => memoryror_202);
    
    memoryrff_166_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya166_Z, B => WriteEnable, Y => 
        memorywre_166);
    
    memory_memory_0_0_sr_RNO_266 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_42, B => memoryro_426, C => 
        memorya426_Z, D => memorya42_Z, Y => memoryror_124);
    
    memoryrff_467 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_467, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_467);
    
    memoryrff_116 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_116, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_116);
    
    memoryrff_82_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya82_Z, B => WriteEnable, Y => 
        memorywre_82);
    
    memory_memory_0_0_sr_RNO_307 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_15, B => memoryro_271, C => 
        memorya271_Z, D => memorya15, Y => memoryror_3);
    
    memoryrff_230 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_230, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_230);
    
    memoryrff_101 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_101, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_101);
    
    memorya268_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya273_4_Z, B => memorya45_3_Z, Y => 
        memorya268_6_Z);
    
    memorya421_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya369_3_Z, B => memorya68_3_Z, Y => 
        memorya421_6_Z);
    
    memory_memory_0_0_sr_RNO_203 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_186, B => memoryro_266, C => 
        memorya266_Z, D => memorya186_Z, Y => memoryror_188);
    
    memoryrff_485 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_485, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_485);
    
    memoryrff_378_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya378_Z, B => WriteEnable, Y => 
        memorywre_378);
    
    memoryrff_103_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya103_Z, B => WriteEnable, Y => 
        memorywre_103);
    
    memory_memory_0_0_sr_RNO_113 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_501, B => memoryro_197, C => 
        memorya501_Z, D => memorya197_Z, Y => memoryror_235);
    
    memoryrff_19 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_19, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_19);
    
    memory_memory_0_0_sr_RNO_55 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_82, B => memoryror_83, C => 
        memoryror_81, D => memoryror_80, Y => memoryror_404);
    
    memoryrff_293_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya305_2_Z, B => WriteEnable, C => 
        memorya292_6_Z, D => memorya261_0_Z, Y => memorywre_293);
    
    memoryrff_305_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya305_Z, B => WriteEnable, Y => 
        memorywre_305);
    
    memorya355 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya116_2_Z, B => memorya355_6_Z, C => 
        InternalAddr2Memory(7), D => memorya379_1_Z, Y => 
        memorya355_Z);
    
    memoryrff_65_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya65_Z, B => WriteEnable, Y => 
        memorywre_65);
    
    memoryrff_126_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya126_Z, B => WriteEnable, Y => 
        memorywre_126);
    
    memory_memory_0_0_sr_RNO_43 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_145, B => memoryror_147, C => 
        memoryror_146, D => memoryror_144, Y => memoryror_420);
    
    memoryrff_406 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_406, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_406);
    
    memorya480 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(4), B => memorya116_2_Z, 
        C => memorya368_6_Z, D => memorya498_3_Z, Y => 
        memorya480_Z);
    
    memorya345 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya86_2_Z, B => memorya345_6_Z, C => 
        InternalAddr2Memory(7), D => memorya121_1_Z, Y => 
        memorya345_Z);
    
    memoryrff_162 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_162, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_162);
    
    memoryrff_432 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_432, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_432);
    
    memoryrff_395 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_395, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_395);
    
    memorya26 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya25_3_Z, B => memorya362_1_Z, C => 
        memorya52_4, D => memorya16_0_Z, Y => memorya26_Z);
    
    memoryrff_434 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_434, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_434);
    
    memorya23 : CFG3
      generic map(INIT => x"20")

      port map(A => memorya20_6_Z, B => InternalAddr2Memory(8), C
         => memorya503_5_Z, Y => memorya23_Z);
    
    memory_memory_0_0_sr_RNO_85 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_217, B => memoryro_473, C => 
        memorya473_Z, D => memorya217_Z, Y => memoryror_221);
    
    memoryrff_5_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya117_1_Z, C => 
        memorya5_0_Z, D => memorya4_6_Z, Y => memorywre_5);
    
    memorya369 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya368_4_Z, B => InternalAddr2Memory(7), 
        C => memorya369_5_Z, D => memorya369_3_Z, Y => 
        memorya369_Z);
    
    memory_memory_0_0_sr_RNO_353 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya102_1_Z, B => memorya8_0_Z, C => 
        memorya4_6_Z, Y => memorya14);
    
    memoryrff_1_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya1_Z, B => WriteEnable, Y => 
        memorywre_1);
    
    memorya77_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya77_2_Z, B => memorya117_1_Z, Y => 
        memorya77_5_Z);
    
    memory_memory_0_0_sr_RNO_69 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_51, B => memoryror_50, C => 
        memoryror_49, D => memoryror_48, Y => memoryror_396);
    
    memoryrff_51 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_51, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_51);
    
    memoryrff_399 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_399, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_399);
    
    memorya391_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya487_4_Z, B => memorya4_3_Z, Y => 
        memorya391_6_Z);
    
    memorya339 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya86_2_Z, B => memorya339_6_Z, C => 
        InternalAddr2Memory(7), D => memorya379_1_Z, Y => 
        memorya339_Z);
    
    memoryrff_317 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_317, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_317);
    
    memorya100_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya102_4_Z, B => memorya84_3_Z, Y => 
        memorya100_6_Z);
    
    memoryrff_26 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_26, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_26);
    
    memorya325 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya261_0_Z, B => memorya368_2_Z, C => 
        memorya197_6_Z, Y => memorya325_Z);
    
    memory_memory_0_0_sr_RNO_242 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_79, B => memoryro_335, C => 
        memorya335_Z, D => memorya79_Z, Y => memoryror_67);
    
    memoryrff_89 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_89, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_89);
    
    memorya117 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya117_1_Z, B => memorya54_2_Z, C => 
        memorya116_4_Z, D => memorya93_0, Y => memorya117_Z);
    
    memory_memory_0_0_sr_RNO_12 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_407, B => memoryror_406, C => 
        memoryror_405, D => memoryror_404, Y => memoryror_485);
    
    memoryrff_461_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya461_Z, B => WriteEnable, Y => 
        memorywre_461);
    
    memoryrff_332 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_332, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_332);
    
    memoryrff_264 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_264, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_264);
    
    memorya78_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya77_2_Z, B => memorya102_1_Z, Y => 
        memorya78_5_Z);
    
    memoryrff_188 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_188, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_188);
    
    memory_memory_0_0_sr_RNO_66 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_114, B => memoryror_112, C => 
        memoryror_113, D => memoryror_115, Y => memoryror_412);
    
    memoryrff_288_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya288_Z, B => WriteEnable, Y => 
        memorywre_288);
    
    memoryrff_287 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_287, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_287);
    
    memoryrff_340 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_340, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_340);
    
    memorya320_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya4_3_Z, B => memorya368_4_Z, Y => 
        memorya320_6_Z);
    
    memoryrff_336 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_336, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_336);
    
    memoryrff_380_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya380_Z, B => WriteEnable, Y => 
        memorywre_380);
    
    memory_memory_0_0_sr_RNO_339 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_388, B => memoryro_20, C => 
        memorya388_Z, D => memorya20, Y => memoryror_25);
    
    memory_memory_0_0_sr_RNO_370 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya4_6_Z, B => memorya379_1_Z, C => 
        memorya3_0_Z, Y => memorya3);
    
    memorya250 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya54_2_Z, B => memorya362_1_Z, C => 
        memorya482_2_Z, D => memorya10_0_Z, Y => memorya250_Z);
    
    memoryrff_421_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya421_Z, B => WriteEnable, Y => 
        memorywre_421);
    
    memory_memory_0_0_sr_RNO_217 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_84, B => memoryro_452, C => 
        memorya452_Z, D => memorya84_Z, Y => memoryror_89);
    
    memoryrff_437 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_437, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_437);
    
    memorya240 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya54_2_Z, C
         => memorya368_6_Z, D => memorya482_2_Z, Y => 
        memorya240_Z);
    
    memoryrff_405 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_405, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_405);
    
    memoryrff_217_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya217_Z, B => WriteEnable, Y => 
        memorywre_217);
    
    memorya55_0 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(3), Y => memorya55_0_Z);
    
    memorya312 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya280_0_Z, B => memorya305_2_Z, C => 
        memorya68_2_Z, D => memorya312_4_Z, Y => memorya312_Z);
    
    memoryrff_389_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya389_Z, B => WriteEnable, Y => 
        memorywre_389);
    
    memorya77_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(3), Y => memorya77_2_Z);
    
    memory_memory_0_0_sr_RNO_99 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_459, B => memoryro_11, C => 
        memorya459_Z, D => memorya11_Z, Y => memoryror_213);
    
    \memory_memory_0_0_OLDA_RNILMUT[0]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(0), C => 
        memory_memory_0_0_OLDA_Z(0), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(0));
    
    \memory_memory_0_0_OLDA_RNIAMT31[14]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(14), C => 
        memory_memory_0_0_OLDA_Z(14), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(14));
    
    memory_memory_0_0_sr_RNO_334 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_263, B => memoryro_23, C => 
        memorya263_Z, D => memorya23_Z, Y => memoryror_30);
    
    memoryrff_220 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_220, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_220);
    
    memorya103_0 : CFG3
      generic map(INIT => x"04")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(6), C => InternalAddr2Memory(8), Y
         => memorya87_0);
    
    memoryrff_49_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya49_Z, B => WriteEnable, Y => 
        memorywre_49);
    
    memorya461 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya45_3_Z, C
         => memorya77_5_Z, D => memorya498_3_Z, Y => memorya461_Z);
    
    memoryrff_113 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_113, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_113);
    
    memorya419 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_1_Z, B => InternalAddr2Memory(6), 
        C => memorya355_6_Z, D => memorya434_2_Z, Y => 
        memorya419_Z);
    
    memorya313 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya312_4_Z, B => InternalAddr2Memory(7), 
        C => memorya121_5_Z, D => memorya369_3_Z, Y => 
        memorya313_Z);
    
    memorya431 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya463_4_Z, 
        C => memorya434_2_Z, D => memorya463_5_Z, Y => 
        memorya431_Z);
    
    memory_memory_0_0_sr_RNO_336 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_277, B => memoryro_21, C => 
        memorya277_Z, D => memorya21, Y => memoryror_27);
    
    memoryrff_15 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_15, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_15);
    
    memoryrff_46 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_46, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_46);
    
    memorya220 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya29_3_Z, C
         => memorya162_2_Z, D => memorya348_5_Z, Y => 
        memorya220_Z);
    
    memoryrff_132 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_132, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_132);
    
    memoryrff_113_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya113_Z, B => WriteEnable, Y => 
        memorywre_113);
    
    memorya338 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya338_6_Z, B => memorya368_2_Z, C => 
        InternalAddr2Memory(7), D => memorya370_1_Z, Y => 
        memorya338_Z);
    
    memory_memory_0_0_sr_RNO_39 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_167, B => memoryror_166, C => 
        memoryror_165, D => memoryror_164, Y => memoryror_425);
    
    memory_memory_0_0_sr_RNO_192 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_256, B => memoryro_48, C => 
        memorya256_Z, D => memorya48, Y => memoryror_130);
    
    memoryrff_367_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya367_Z, B => WriteEnable, Y => 
        memorywre_367);
    
    memoryrff_17 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_17, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_17);
    
    memory_memory_0_0_sr_RNO_96 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_173, B => memoryro_477, C => 
        memorya477_Z, D => memorya173_Z, Y => memoryror_214);
    
    memoryrff_315_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya315_Z, B => WriteEnable, Y => 
        memorywre_315);
    
    memoryrff_480_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya480_Z, B => WriteEnable, Y => 
        memorywre_480);
    
    memoryrff_265 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_265, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_265);
    
    memory_memory_0_0_sr_RNO_129 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_212, B => memoryro_260, C => 
        memorya260_Z, D => memorya212_Z, Y => memoryror_201);
    
    memoryrff_422 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_422, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_422);
    
    memory_memory_0_0_sr_RNO_40 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_157, B => memoryror_156, C => 
        memoryror_159, D => memoryror_158, Y => memoryror_423);
    
    memory_memory_0_0_sr_RNO_120 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_455, B => memoryro_151, C => 
        memorya455_Z, D => memorya151_Z, Y => memoryror_206);
    
    memoryrff_355 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_355, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_355);
    
    memorya84_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(1), Y => memorya84_3_Z);
    
    memoryrff_182_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya182_Z, B => WriteEnable, Y => 
        memorywre_182);
    
    memoryrff_424 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_424, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_424);
    
    memoryrff_375 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_375, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_375);
    
    memory_memory_0_0_sr_RNO_78 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_47, B => memoryror_45, C => 
        memoryror_46, D => memoryror_44, Y => memoryror_395);
    
    memoryrff_304_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya304_Z, B => WriteEnable, Y => 
        memorywre_304);
    
    memory_memory_0_0_sr_RNO_36 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_168, B => memoryror_171, C => 
        memoryror_170, D => memoryror_169, Y => memoryror_426);
    
    memory_memory_0_0_sr_RNO_162 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_443, B => memoryro_91, C => 
        memorya443_Z, D => memorya91_Z, Y => memoryror_165);
    
    memory_memory_0_0_sr_RNO : CFG4
      generic map(INIT => x"0001")

      port map(A => memoryror_507, B => memoryror_506, C => 
        memoryror_505, D => memoryror_504, Y => memoryror_i);
    
    memorya96 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya368_4_Z, B => memorya102_4_Z, C => 
        memorya116_2_Z, D => memorya20_0_Z, Y => memorya96_Z);
    
    memorya178 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya370_1_Z, B => InternalAddr2Memory(8), 
        C => memorya306_6_Z, D => memorya434_2_Z, Y => 
        memorya178_Z);
    
    memory_memory_0_0_sr_RNO_350 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya167_3_Z, B => memorya199_0_Z, C => 
        memorya455_5_Z, Y => memorya199);
    
    memoryrff_455_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya455_Z, B => WriteEnable, Y => 
        memorywre_455);
    
    memoryrff_42_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya42_Z, B => WriteEnable, Y => 
        memorywre_42);
    
    memoryrff_23 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_23, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_23);
    
    memoryrff_108 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_108, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_108);
    
    memoryrff_435_RNO : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya499_5_Z, B => memorya435_6_Z, C => 
        InternalAddr2Memory(6), D => WriteEnable, Y => 
        memorywre_435);
    
    memoryrff_359 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_359, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_359);
    
    memorya93 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya117_1_Z, B => memorya125_2_Z, C => 
        memorya93_0, D => memorya68_4_Z, Y => memorya93_Z);
    
    memorya481_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya482_2_Z, B => memorya353_1_Z, Y => 
        memorya481_5_Z);
    
    memoryrff_327_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya327_Z, B => WriteEnable, Y => 
        memorywre_327);
    
    memoryrff_234 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_234, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_234);
    
    memoryrff_61_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya61_Z, B => WriteEnable, Y => 
        memorywre_61);
    
    memoryrff_379 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_379, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_379);
    
    memoryrff_207 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_207, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_207);
    
    memoryrff_85 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_85, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_85);
    
    memory_memory_0_0_sr_RNO_378 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya464_0_Z, B => memorya368_6_Z, Y => 
        memorya464);
    
    memorya67 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya67_2_Z, B => memorya68_6_Z, C => 
        InternalAddr2Memory(8), D => memorya379_1_Z, Y => 
        memorya67_Z);
    
    memory_memory_0_0_sr_RNO_244 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_408, B => memoryro_24, C => 
        memorya408_Z, D => memorya24_Z, Y => memoryror_111);
    
    memoryrff_322 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_322, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_322);
    
    memoryrff_87 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_87, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_87);
    
    memoryrff_7 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_7, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_7);
    
    memoryrff_384 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_384, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_384);
    
    \memory_memory_0_0_OLDA[29]\ : SLE
      port map(D => \InternalDataFromMem\(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(29));
    
    memoryrff_504_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya504_Z, B => WriteEnable, Y => 
        memorywre_504);
    
    memoryrff_467_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya467_Z, B => WriteEnable, Y => 
        memorywre_467);
    
    memory_memory_0_0_sr_RNO_145 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_244, B => memoryro_308, C => 
        memorya308_Z, D => memorya244_Z, Y => memoryror_249);
    
    memorya473 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya86_2_Z, B => memorya441_6_Z, C => 
        InternalAddr2Memory(5), D => memorya121_1_Z, Y => 
        memorya473_Z);
    
    memorya45_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(3), Y => memorya45_2_Z);
    
    memorya172 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya68_2_Z, C
         => memorya289_4_Z, D => memorya428_5_Z, Y => 
        memorya172_Z);
    
    memory_memory_0_0_sr_RNO_345 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya264_6_Z, B => memorya395_2_Z, C => 
        memorya20_0_Z, Y => memorya136);
    
    memory_memory_0_0_sr_RNO_241 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_418, B => memoryro_194, C => 
        memorya418_Z, D => memorya194_Z, Y => memoryror_64);
    
    memoryrff_326 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_326, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_326);
    
    memorya368_0 : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory(7), B => memorya54_2_Z, C
         => memorya368_2_Z, Y => memorya368_0_Z);
    
    memorya188 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya316_4_Z, 
        C => memorya162_2_Z, D => memorya380_5_Z, Y => 
        memorya188_Z);
    
    memory_memory_0_0_sr : SLE
      port map(D => memoryror_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => memory_memory_0_0_sr_Z);
    
    memory_memory_0_0_sr_RNO_321 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_420, B => memoryro_36, C => 
        memorya420_Z, D => memorya36, Y => memoryror_41);
    
    memoryrff_170_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya170_Z, B => WriteEnable, Y => 
        memorywre_170);
    
    memorya264_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya273_4_Z, B => memorya41_3_Z, Y => 
        memorya264_6_Z);
    
    memory_memory_0_0_sr_RNO_240 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_416, B => memoryro_240, C => 
        memorya416_Z, D => memorya240_Z, Y => memoryror_66);
    
    memoryrff_427 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_427, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_427);
    
    memory_memory_0_0_sr_RNO_309 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_301, B => memoryro_29, C => 
        memorya301_Z, D => memorya29_Z, Y => memoryror_38);
    
    memory_memory_0_0_sr_RNO_286 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_317, B => memoryro_13, C => 
        memorya317_Z, D => memorya13_Z, Y => memoryror_54);
    
    memoryrff_427_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya427_Z, B => WriteEnable, Y => 
        memorywre_427);
    
    memorya510 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya116_2_Z, B => InternalAddr2Memory(0), 
        C => memorya126_5_Z, D => memorya498_3_Z, Y => 
        memorya510_Z);
    
    memory_memory_0_0_sr_RNO_298 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_261, B => memoryro_5, C => 
        memorya261_Z, D => memorya5, Y => memoryror_11);
    
    memoryrff_368_RNO : CFG3
      generic map(INIT => x"80")

      port map(A => WriteEnable, B => memorya368_6_Z, C => 
        memorya368_0_Z, Y => memorywre_368);
    
    memorya68 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya68_4_Z, B => memorya20_0_Z, C => 
        memorya68_3_Z, D => memorya68_1_Z, Y => memorya68_Z);
    
    memoryrff_88_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya88_Z, B => WriteEnable, Y => 
        memorywre_88);
    
    memoryrff_20_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya116_1_Z, B => WriteEnable, C => 
        memorya20_0_Z, D => memorya20_6_Z, Y => memorywre_20);
    
    memoryrff_119 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_119, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_119);
    
    memorya277 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya273_4_Z, B => memorya84_3_Z, C => 
        memorya261_0_Z, D => memorya278_2_Z, Y => memorya277_Z);
    
    memorya268 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya268_6_Z, B => memorya268_0_Z, C => 
        memorya370_3_Z, Y => memorya268_Z);
    
    memoryrff_483_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya483_Z, B => WriteEnable, Y => 
        memorywre_483);
    
    memory_memory_0_0_sr_RNO_51 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_186, B => memoryror_184, C => 
        memoryror_185, D => memoryror_187, Y => memoryror_430);
    
    memorya238 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya46_3_Z, C
         => memorya110_5_Z, D => memorya482_2_Z, Y => 
        memorya238_Z);
    
    memorya9_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya121_1_Z, B => InternalAddr2Memory(8), 
        Y => memorya9_0_Z);
    
    memorya262 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_1_Z, B => InternalAddr2Memory(7), 
        C => memorya257_6_Z, D => memorya370_3_Z, Y => 
        memorya262_Z);
    
    memorya162_2 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(0), Y => memorya162_2_Z);
    
    memoryrff_479_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya479_Z, B => WriteEnable, Y => 
        memorywre_479);
    
    memoryrff_290 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_290, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_290);
    
    memorya232 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya45_2_Z, C
         => memorya360_6_Z, D => memorya482_2_Z, Y => 
        memorya232_Z);
    
    memoryrff_87_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya87_Z, B => WriteEnable, Y => 
        memorywre_87);
    
    memoryrff_43 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_43, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_43);
    
    memorya202_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya4_3_Z, B => memorya354_3_Z, Y => 
        memorya202_6_Z);
    
    memorya483 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(4), B => memorya379_1_Z, 
        C => memorya116_2_Z, D => memorya435_6_Z, Y => 
        memorya483_Z);
    
    memory_memory_0_0_sr_RNO_304 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_176, B => memoryro_448, C => 
        memorya448_Z, D => memorya176_Z, Y => memoryror_2);
    
    memorya253 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya125_2_Z, B => memorya117_1_Z, C => 
        memorya193_2_Z, D => memorya111_0_Z, Y => memorya253_Z);
    
    memorya182 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya162_2_Z, B => memorya118_5_Z, C => 
        InternalAddr2Memory(8), D => memorya304_4_Z, Y => 
        memorya182_Z);
    
    memory_memory_0_0_sr_RNO_268 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_384, B => memoryro_192, C => 
        memorya384_Z, D => memorya192_Z, Y => memoryror_114);
    
    memorya377 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya57_3_Z, B => InternalAddr2Memory(7), C
         => memorya121_5_Z, D => memorya368_2_Z, Y => 
        memorya377_Z);
    
    memory_memory_0_0_sr_RNO_358 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya362_1_Z, B => memorya10_0_Z, C => 
        memorya4_6_Z, Y => memorya10);
    
    \memory_memory_0_0_OLDA[27]\ : SLE
      port map(D => \InternalDataFromMem\(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(27));
    
    memorya243 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya3_0_Z, B => memorya482_2_Z, C => 
        memorya499_5_Z, Y => memorya243_Z);
    
    memorya490 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(4), B => memorya362_1_Z, 
        C => memorya116_2_Z, D => memorya498_6_Z, Y => 
        memorya490_Z);
    
    memoryrff_235 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_235, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_235);
    
    memoryrff_122 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_122, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_122);
    
    memorya204 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya364_1_Z, 
        C => memorya204_6_Z, D => memorya482_2_Z, Y => 
        memorya204_Z);
    
    memoryrff_328_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya328_Z, B => WriteEnable, Y => 
        memorywre_328);
    
    memory_memory_0_0_sr_RNO_306 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_481, B => memoryro_65, C => 
        memorya481_Z, D => memorya65_Z, Y => memoryror_1);
    
    memory_memory_0_0_sr_RNO_81 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_21, B => memoryror_22, C => 
        memoryror_20, D => memoryror_23, Y => memoryror_389);
    
    memory_memory_0_0_sr_RNO_174 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_275, B => memoryro_147, C => 
        memorya275_Z, D => memorya147_Z, Y => memoryror_152);
    
    memorya370_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya370_3_Z, B => memorya368_4_Z, Y => 
        memorya370_6_Z);
    
    memory_memory_0_0_sr_RNO_313 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_480, B => memoryro_144, C => 
        memorya480_Z, D => memorya144, Y => memoryror_34);
    
    memoryrff_368 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_368, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_368);
    
    memoryrff_50_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya50_Z, B => WriteEnable, Y => 
        memorywre_50);
    
    memoryrff_107_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya107_Z, B => WriteEnable, Y => 
        memorywre_107);
    
    memoryrff_492 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_492, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_492);
    
    memoryrff_14 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_14, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_14);
    
    memorya287 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya273_4_Z, 
        C => memorya278_2_Z, D => memorya463_5_Z, Y => 
        memorya287_Z);
    
    memoryrff_304 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_304, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_304);
    
    memoryrff_179_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya179_Z, B => WriteEnable, Y => 
        memorywre_179);
    
    memoryrff_180 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_180, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_180);
    
    memoryrff_494 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_494, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_494);
    
    memorya405 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya20_3_Z, B => InternalAddr2Memory(6), C
         => memorya149_5_Z, D => memorya369_3_Z, Y => 
        memorya405_Z);
    
    memoryrff_22 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_22, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_22);
    
    memory_memory_0_0_sr_RNO_147 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_438, B => memoryro_246, C => 
        memorya438_Z, D => memorya246_Z, Y => memoryror_250);
    
    memoryrff_314_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya314_Z, B => WriteEnable, Y => 
        memorywre_314);
    
    memorya223 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya223_0_Z, 
        C => memorya86_2_Z, D => memorya463_5_Z, Y => 
        memorya223_Z);
    
    \memory_memory_0_0_OLDA[21]\ : SLE
      port map(D => \InternalDataFromMem\(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(21));
    
    memoryrff_442_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya442_Z, B => WriteEnable, Y => 
        memorywre_442);
    
    memoryrff_224 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_224, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_224);
    
    memoryrff_209_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya209_Z, B => WriteEnable, Y => 
        memorywre_209);
    
    memory_memory_0_0_sr_RNO_293 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_9, B => memoryro_265, C => 
        memorya265_Z, D => memorya9, Y => memoryror_13);
    
    memoryrff_345 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_345, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_345);
    
    memorya387 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_1_Z, B => InternalAddr2Memory(6), 
        C => memorya320_6_Z, D => memorya498_3_Z, Y => 
        memorya387_Z);
    
    memoryrff_419 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_419, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_419);
    
    memorya315 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya312_4_Z, 
        C => memorya305_2_Z, D => memorya315_5_Z, Y => 
        memorya315_Z);
    
    memory_memory_0_0_sr_RNO_367 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya199_0_Z, B => memorya331_5_Z, C => 
        memorya211_3_Z, Y => memorya203);
    
    memoryrff_392 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_392, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_392);
    
    memory_memory_0_0_sr_RNO_68 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_60, B => memoryror_61, C => 
        memoryror_63, D => memoryror_62, Y => memoryror_399);
    
    memoryrff_468 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_468, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_468);
    
    memoryrff_349 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_349, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_349);
    
    memory_memory_0_0_sr_RNO_263 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_139, B => memoryro_267, C => 
        memorya267_Z, D => memorya139_Z, Y => memoryror_117);
    
    memoryrff_84 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_84, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_84);
    
    memorya47 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya47_0_Z, C
         => memorya463_5_Z, D => memorya52_4, Y => memorya47_Z);
    
    memorya371 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya368_4_Z, 
        C => memorya368_2_Z, D => memorya499_5_Z, Y => 
        memorya371_Z);
    
    memoryrff_396 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_396, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_396);
    
    memory_memory_0_0_sr_RNO_154 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_288, B => memoryro_16, C => 
        memorya288_Z, D => memorya16, Y => memoryror_162);
    
    memoryrff_488_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya488_Z, B => WriteEnable, Y => 
        memorywre_488);
    
    memorya11 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya11_0_Z, B => InternalAddr2Memory(8), C
         => memorya379_1_Z, D => memorya4_6_Z, Y => memorya11_Z);
    
    memoryrff_497 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_497, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_497);
    
    memoryrff_257_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya257_Z, B => WriteEnable, Y => 
        memorywre_257);
    
    memoryrff_237_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya237_Z, B => WriteEnable, Y => 
        memorywre_237);
    
    memorya83_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya68_4_Z, B => memorya368_4_Z, Y => 
        memorya83_6_Z);
    
    memorya379_4 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(2), Y => memorya379_4_Z);
    
    memoryrff_492_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya492_Z, B => WriteEnable, Y => 
        memorywre_492);
    
    memoryrff_281_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya281_Z, B => WriteEnable, Y => 
        memorywre_281);
    
    memorya271 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya463_4_Z, 
        C => memorya273_4_Z, D => memorya463_5_Z, Y => 
        memorya271_Z);
    
    memory_memory_0_0_sr_RNO_222 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_93, B => memoryro_349, C => 
        memorya349_Z, D => memorya93_Z, Y => memoryror_86);
    
    memoryrff_250 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_250, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_250);
    
    memoryrff_42 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_42, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_42);
    
    memoryrff_270 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_270, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_270);
    
    memoryrff_200_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya200_Z, B => WriteEnable, Y => 
        memorywre_200);
    
    memoryrff_383_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya383_Z, B => WriteEnable, Y => 
        memorywre_383);
    
    memory_memory_0_0_sr_RNO_98 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_284, B => memoryro_204, C => 
        memorya284_Z, D => memorya204_Z, Y => memoryror_212);
    
    memoryrff_100 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_100, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_100);
    
    memorya381 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya116_2_Z, 
        C => memorya369_3_Z, D => memorya381_5_Z, Y => 
        memorya381_Z);
    
    memorya254 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya116_2_Z, B => InternalAddr2Memory(8), 
        C => memorya126_5_Z, D => memorya162_2_Z, Y => 
        memorya254_Z);
    
    \memory_memory_0_0_OLDA[2]\ : SLE
      port map(D => \InternalDataFromMem\(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(2));
    
    memoryrff_338 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_338, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_338);
    
    memoryrff_225 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_225, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_225);
    
    memorya210 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya370_1_Z, 
        C => memorya338_6_Z, D => memorya482_2_Z, Y => 
        memorya210_Z);
    
    memoryrff_73_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya73_Z, B => WriteEnable, Y => 
        memorywre_73);
    
    memoryrff_192 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_192, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_192);
    
    memoryrff_153_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya153_Z, B => WriteEnable, Y => 
        memorywre_153);
    
    memorya244 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya5_0_Z, B => memorya116_1_Z, C => 
        memorya162_2_Z, D => memorya116_2_Z, Y => memorya244_Z);
    
    memoryrff_133_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya133_Z, B => WriteEnable, Y => 
        memorywre_133);
    
    memorya111_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya116_2_Z, B => InternalAddr2Memory(8), 
        Y => memorya111_0_Z);
    
    memory_memory_0_0_sr_RNO_310 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_347, B => memoryro_219, C => 
        memorya347_Z, D => memorya219_Z, Y => memoryror_37);
    
    memoryrff_0_RNO : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya368_6_Z, B => memorya4_6_Z, C => 
        InternalAddr2Memory(8), D => WriteEnable, Y => 
        memorywre_0);
    
    memoryrff_355_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya355_Z, B => WriteEnable, Y => 
        memorywre_355);
    
    memoryrff_452 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_452, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_452);
    
    memoryrff_335_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya335_Z, B => WriteEnable, Y => 
        memorywre_335);
    
    memory_memory_0_0_sr_RNO_141 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_446, B => memoryro_126, C => 
        memorya446_Z, D => memorya126_Z, Y => memoryror_247);
    
    memoryrff_346_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya346_Z, B => WriteEnable, Y => 
        memorywre_346);
    
    memory_memory_0_0_sr_RNO_38 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_174, B => memoryror_173, C => 
        memoryror_175, D => memoryror_172, Y => memoryror_427);
    
    memory_memory_0_0_sr_RNO_182 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_131, B => memoryro_259, C => 
        memorya259_Z, D => memorya131_Z, Y => memoryror_136);
    
    memoryrff_48_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya54_2_Z, B => WriteEnable, C => 
        memorya51_6_Z, D => memorya20_0_Z, Y => memorywre_48);
    
    memoryrff_472 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_472, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_472);
    
    memoryrff_117_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya117_Z, B => WriteEnable, Y => 
        memorywre_117);
    
    memorya281 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya121_1_Z, 
        C => memorya278_2_Z, D => memorya280_6_Z, Y => 
        memorya281_Z);
    
    memoryrff_454 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_454, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_454);
    
    memorya455 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya68_3_Z, C
         => memorya455_5_Z, D => memorya498_3_Z, Y => 
        memorya455_Z);
    
    memorya380_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya54_2_Z, B => memorya364_1_Z, Y => 
        memorya380_5_Z);
    
    memory_memory_0_0_sr_RNO_136 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_376, B => memoryro_136, C => 
        memorya376_Z, D => memorya136, Y => memoryror_255);
    
    memorya46_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(0), Y => memorya46_3_Z);
    
    memory_memory_0_0_sr_RNO_27 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_233, B => memoryror_235, C => 
        memoryror_234, D => memoryror_232, Y => memoryror_442);
    
    memoryrff_474 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_474, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_474);
    
    memoryrff_188_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya188_Z, B => WriteEnable, Y => 
        memorywre_188);
    
    memorya445 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya369_3_Z, B => memorya381_5_Z, C => 
        InternalAddr2Memory(6), D => memorya434_2_Z, Y => 
        memorya445_Z);
    
    memoryrff_29 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_29, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_29);
    
    memoryrff_47_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya47_Z, B => WriteEnable, Y => 
        memorywre_47);
    
    memoryrff_294 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_294, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_294);
    
    memorya273_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(5), Y => memorya273_4_Z);
    
    memorya224 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya116_2_Z, 
        C => memorya162_2_Z, D => memorya353_6_Z, Y => 
        memorya224_Z);
    
    memorya477 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya369_3_Z, 
        C => memorya381_5_Z, D => memorya482_2_Z, Y => 
        memorya477_Z);
    
    memoryrff_438 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_438, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_438);
    
    memoryrff_219_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya219_Z, B => WriteEnable, Y => 
        memorywre_219);
    
    memoryrff_203_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya211_3_Z, B => WriteEnable, C => 
        memorya331_5_Z, D => memorya199_0_Z, Y => memorywre_203);
    
    memorya5_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya84_3_Z, B => InternalAddr2Memory(8), Y
         => memorya5_0_Z);
    
    memorya33 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya57_3_Z, B => memorya36_6_Z, C => 
        InternalAddr2Memory(8), D => memorya353_1_Z, Y => 
        memorya33_Z);
    
    memoryrff_352 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_352, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_352);
    
    memoryrff_372 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_372, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_372);
    
    memoryrff_160_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya160_Z, B => WriteEnable, Y => 
        memorywre_160);
    
    memorya176 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya304_4_Z, B => memorya57_3_Z, C => 
        memorya63_0, D => memorya162_2_Z, Y => memorya176_Z);
    
    memorya499_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya54_2_Z, B => memorya379_1_Z, Y => 
        memorya499_5_Z);
    
    memory_memory_0_0_sr_RNO_49 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_191, B => memoryror_190, C => 
        memoryror_189, D => memoryror_188, Y => memoryror_431);
    
    memorya101 : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory(8), B => memorya100_6_Z, 
        C => memorya101_5_Z, Y => memorya101_Z);
    
    memorya198 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya102_1_Z, 
        C => memorya326_6_Z, D => memorya482_2_Z, Y => 
        memorya198_Z);
    
    memorya425 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya121_1_Z, B => InternalAddr2Memory(6), 
        C => memorya361_6_Z, D => memorya434_2_Z, Y => 
        memorya425_Z);
    
    memorya312_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(2), Y => memorya312_4_Z);
    
    memorya126_0 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(0), Y => memorya126_0_Z);
    
    memoryrff_356 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_356, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_356);
    
    memorya170 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya362_1_Z, B => InternalAddr2Memory(8), 
        C => memorya298_6_Z, D => memorya434_2_Z, Y => 
        memorya170_Z);
    
    memory_memory_0_0_sr_RNO_138 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_167, B => memoryro_503, C => 
        memorya503_Z, D => memorya167_Z, Y => memoryror_254);
    
    memorya504 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(2), B => memorya125_2_Z, 
        C => memorya116_2_Z, D => memorya504_6_Z, Y => 
        memorya504_Z);
    
    memoryrff_396_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya396_Z, B => WriteEnable, Y => 
        memorywre_396);
    
    memoryrff_376 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_376, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_376);
    
    memoryrff_469_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya469_Z, B => WriteEnable, Y => 
        memorywre_469);
    
    memorya69 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya117_1_Z, B => InternalAddr2Memory(8), 
        C => memorya68_6_Z, D => memorya117_3_Z, Y => memorya69_Z);
    
    \memory_memory_0_0_OLDA[7]\ : SLE
      port map(D => \InternalDataFromMem\(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(7));
    
    memoryrff_457 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_457, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_457);
    
    memory_memory_0_0_sr_RNO_46 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_140, B => memoryror_143, C => 
        memoryror_142, D => memoryror_141, Y => memoryror_419);
    
    memorya487 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya487_4_Z, B => InternalAddr2Memory(4), 
        C => memorya482_2_Z, D => memorya487_5_Z, Y => 
        memorya487_Z);
    
    memoryrff_120_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya120_Z, B => WriteEnable, Y => 
        memorywre_120);
    
    memorya300 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya68_2_Z, B => memorya289_4_Z, C => 
        memorya268_0_Z, D => memorya305_2_Z, Y => memorya300_Z);
    
    \memory_memory_0_0_OLDA[5]\ : SLE
      port map(D => \InternalDataFromMem\(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(5));
    
    memoryrff_477 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_477, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_477);
    
    memoryrff_481 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_481, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_481);
    
    memoryrff_269 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_269, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_269);
    
    memory_memory_0_0_sr_RNO_318 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_55, B => memoryro_311, C => 
        memorya311_Z, D => memorya55_Z, Y => memoryror_46);
    
    memoryrff_486_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya486_Z, B => WriteEnable, Y => 
        memorywre_486);
    
    memoryrff_9 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_9, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_9);
    
    memorya493 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(4), B => memorya369_3_Z, 
        C => memorya45_5_Z, D => memorya482_2_Z, Y => 
        memorya493_Z);
    
    memorya186 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya312_4_Z, 
        C => memorya162_2_Z, D => memorya378_5_Z, Y => 
        memorya186_Z);
    
    memory_memory_0_0_sr_RNO_342 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya227_0_Z, B => memorya101_5_Z, C => 
        memorya193_2_Z, Y => memorya229);
    
    memory_memory_0_0_sr_RNO_224 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_224, B => memoryro_432, C => 
        memorya432, D => memorya224_Z, Y => memoryror_82);
    
    memoryrff_281 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_281, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_281);
    
    memorya192 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_2_Z, B => InternalAddr2Memory(8), C
         => memorya320_6_Z, D => memorya482_2_Z, Y => 
        memorya192_Z);
    
    memory_memory_0_0_sr_RNO_25 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_230, B => memoryror_229, C => 
        memoryror_228, D => memoryror_231, Y => memoryror_441);
    
    memoryrff_382_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya382_Z, B => WriteEnable, Y => 
        memorywre_382);
    
    memorya462 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya46_3_Z, B => InternalAddr2Memory(5), C
         => memorya78_5_Z, D => memorya498_3_Z, Y => memorya462_Z);
    
    memory_memory_0_0_sr_RNO_288 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_310, B => memoryro_54, C => 
        memorya310_Z, D => memorya54_Z, Y => memoryror_58);
    
    memoryrff_475_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya475_Z, B => WriteEnable, Y => 
        memorywre_475);
    
    memoryrff_49 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_49, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_49);
    
    memoryrff_429_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya429_Z, B => WriteEnable, Y => 
        memorywre_429);
    
    memoryrff_210_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya210_Z, B => WriteEnable, Y => 
        memorywre_210);
    
    memoryrff_166 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_166, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_166);
    
    memorya180 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya68_2_Z, C
         => memorya304_4_Z, D => memorya436_5_Z, Y => 
        memorya180_Z);
    
    memoryrff_169_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya169_Z, B => WriteEnable, Y => 
        memorywre_169);
    
    memory_memory_0_0_sr_RNO_125 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_66, B => memoryro_258, C => 
        memorya258_Z, D => memorya66_Z, Y => memoryror_192);
    
    memoryrff_328 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_328, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_328);
    
    memoryrff_152 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_152, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_152);
    
    memory_memory_0_0_sr_RNO_325 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_160, B => memoryro_464, C => 
        memorya464, D => memorya160_Z, Y => memoryror_18);
    
    \memory_memory_0_0_OLDA[13]\ : SLE
      port map(D => \InternalDataFromMem\(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(13));
    
    memory_memory_0_0_sr_RNO_221 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_60, B => memoryro_476, C => 
        memorya476_Z, D => memorya60_Z, Y => memoryror_84);
    
    memory_memory_0_0_sr_RNO_0 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_493, B => memoryror_494, C => 
        memoryror_492, D => memoryror_495, Y => memoryror_507);
    
    memoryrff_295 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_295, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_295);
    
    memoryrff_240 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_240, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_240);
    
    memoryrff_172 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_172, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_172);
    
    memorya366 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya46_3_Z, B => InternalAddr2Memory(7), C
         => memorya110_5_Z, D => memorya368_2_Z, Y => 
        memorya366_Z);
    
    memorya297 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya121_1_Z, B => InternalAddr2Memory(7), 
        C => memorya296_6_Z, D => memorya305_2_Z, Y => 
        memorya297_Z);
    
    memoryrff_74_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya74_Z, B => WriteEnable, Y => 
        memorywre_74);
    
    memorya76 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya84_2_Z, B => memorya45_3_Z, C => 
        memorya12_0_Z, D => memorya68_4_Z, Y => memorya76_Z);
    
    memorya408 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya125_2_Z, 
        C => memorya344_6_Z, D => memorya498_3_Z, Y => 
        memorya408_Z);
    
    memorya336 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya86_2_Z, C
         => memorya336_6_Z, D => memorya370_3_Z, Y => 
        memorya336_Z);
    
    memorya304 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya54_2_Z, B => InternalAddr2Memory(7), C
         => memorya304_6_Z, D => memorya370_3_Z, Y => 
        memorya304_Z);
    
    memory_memory_0_0_sr_RNO_220 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_350, B => memoryro_222, C => 
        memorya350_Z, D => memorya222_Z, Y => memoryror_87);
    
    memorya73 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya117_3_Z, B => memorya41_3_Z, C => 
        memorya9_0_Z, D => memorya68_4_Z, Y => memorya73_Z);
    
    GND_Z : GND
      port map(Y => \GND\);
    
    memoryrff_25 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_25, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_25);
    
    memoryrff_129_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya129_Z, B => WriteEnable, Y => 
        memorywre_129);
    
    memorya397 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya117_1_Z, B => InternalAddr2Memory(6), 
        C => memorya333_6_Z, D => memorya395_2_Z, Y => 
        memorya397_Z);
    
    memorya265 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya121_1_Z, B => InternalAddr2Memory(7), 
        C => memorya264_6_Z, D => memorya369_3_Z, Y => 
        memorya265_Z);
    
    memory_memory_0_0_sr_RNO_13 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_401, B => memoryror_402, C => 
        memoryror_403, D => memoryror_400, Y => memoryror_484);
    
    memorya235 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya233_0_Z, B => memorya299_5_Z, C => 
        memorya482_2_Z, Y => memorya235_Z);
    
    memorya213 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya86_2_Z, B => memorya117_1_Z, C => 
        memorya211_0_Z, D => memorya193_2_Z, Y => memorya213_Z);
    
    memory_memory_0_0_sr_RNO_369 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya117_1_Z, B => memorya5_0_Z, C => 
        memorya4_6_Z, Y => memorya5);
    
    memoryrff_71 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_71, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_71);
    
    memoryrff_354_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya354_Z, B => WriteEnable, Y => 
        memorywre_354);
    
    memoryrff_254 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_254, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_254);
    
    memoryrff_442 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_442, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_442);
    
    memoryrff_334_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya334_Z, B => WriteEnable, Y => 
        memorywre_334);
    
    memoryrff_27 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_27, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_27);
    
    memorya105 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya116_2_Z, B => memorya105_6_Z, C => 
        InternalAddr2Memory(8), D => memorya121_1_Z, Y => 
        memorya105_Z);
    
    memory_memory_0_0_sr_RNO_106 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_236, B => memoryro_300, C => 
        memorya300_Z, D => memorya236_Z, Y => memoryror_228);
    
    memoryrff_428 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_428, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_428);
    
    memoryrff_274 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_274, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_274);
    
    memoryrff_60_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya60_Z, B => WriteEnable, Y => 
        memorywre_60);
    
    memoryrff_444 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_444, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_444);
    
    memoryrff_248_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya248_Z, B => WriteEnable, Y => 
        memorywre_248);
    
    memoryrff_213_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya213_Z, B => WriteEnable, Y => 
        memorywre_213);
    
    memoryrff_56 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_56, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_56);
    
    memoryrff_213 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_213, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_213);
    
    memorya163 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_1_Z, B => InternalAddr2Memory(8), 
        C => memorya289_6_Z, D => memorya434_2_Z, Y => 
        memorya163_Z);
    
    memoryrff_367 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_367, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_367);
    
    memoryrff_340_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya340_Z, B => WriteEnable, Y => 
        memorywre_340);
    
    memoryrff_13_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya13_Z, B => WriteEnable, Y => 
        memorywre_13);
    
    memorya116_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(4), B => 
        InternalAddr2Memory(2), Y => memorya116_1_Z);
    
    memory_memory_0_0_sr_RNO_283 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_178, B => memoryro_498, C => 
        memorya498_Z, D => memorya178_Z, Y => memoryror_48);
    
    memorya133 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya117_1_Z, 
        C => memorya193_2_Z, D => memorya257_6_Z, Y => 
        memorya133_Z);
    
    memorya151 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya167_3_Z, 
        C => memorya273_4_Z, D => memorya503_5_Z, Y => 
        memorya151_Z);
    
    memory_memory_0_0_sr_RNO_364 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya57_3_Z, B => memorya8_0_Z, C => 
        memorya4_6_Z, Y => memorya8);
    
    memory_memory_0_0_sr_RNO_114 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_230, B => memoryro_422, C => 
        memorya422_Z, D => memorya230, Y => memoryror_234);
    
    memorya141 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya117_1_Z, B => InternalAddr2Memory(8), 
        C => memorya268_6_Z, D => memorya395_2_Z, Y => 
        memorya141_Z);
    
    memoryrff_401 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_401, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_401);
    
    memoryrff_381_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya381_Z, B => WriteEnable, Y => 
        memorywre_381);
    
    memoryrff_342 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_342, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_342);
    
    memorya278_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya273_4_Z, B => memorya102_3_Z, Y => 
        memorya278_6_Z);
    
    memory_memory_0_0_sr_RNO_366 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya68_3_Z, B => memorya273_4_Z, C => 
        memorya128_0_Z, Y => memorya128);
    
    memoryrff_349_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya349_Z, B => WriteEnable, Y => 
        memorywre_349);
    
    memoryrff_201 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_201, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_201);
    
    memorya361_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya369_3_Z, B => memorya41_3_Z, Y => 
        memorya361_6_Z);
    
    memorya2_0 : CFG2
      generic map(INIT => x"4")

      port map(A => InternalAddr2Memory(0), B => 
        InternalAddr2Memory(1), Y => memorya2_0_Z);
    
    memorya1 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya1_0_Z, B => InternalAddr2Memory(8), C
         => memorya368_4_Z, D => memorya4_6_Z, Y => memorya1_Z);
    
    memoryrff_4_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya4_Z, B => WriteEnable, Y => 
        memorywre_4);
    
    memoryrff_239 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_239, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_239);
    
    memory_memory_0_0_sr_RNO_127 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_321, B => memoryro_193, C => 
        memorya321_Z, D => memorya193_Z, Y => memoryror_193);
    
    memory_memory_0_0_sr_RNO_108 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_487, B => memoryro_183, C => 
        memorya487_Z, D => memorya183_Z, Y => memoryror_238);
    
    memorya350 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya30_3_Z, B => InternalAddr2Memory(7), C
         => memorya126_5_Z, D => memorya368_2_Z, Y => 
        memorya350_Z);
    
    memoryrff_380 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_380, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_380);
    
    memorya434_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(5), Y => memorya434_2_Z);
    
    memorya340 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya276_0_Z, B => memorya340_6_Z, C => 
        memorya368_2_Z, Y => memorya340_Z);
    
    memoryrff_346 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_346, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_346);
    
    memory_memory_0_0_sr_RNO_249 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_100, B => memoryro_484, C => 
        memorya484_Z, D => memorya100_Z, Y => memoryror_105);
    
    memory_memory_0_0_sr_RNO_245 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_103, B => memoryro_359, C => 
        memorya359_Z, D => memorya103_Z, Y => memoryror_110);
    
    \memory_memory_0_0_OLDA_RNIQRUT[5]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(5), C => 
        memory_memory_0_0_OLDA_Z(5), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(5));
    
    memorya121 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya121_1_Z, B => memorya54_2_Z, C => 
        memorya121_4_Z, D => memorya93_0, Y => memorya121_Z);
    
    memoryrff_505_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya505_Z, B => WriteEnable, Y => 
        memorywre_505);
    
    memorya66_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(1), Y => memorya66_1_Z);
    
    \memory_memory_0_0_OLDA[6]\ : SLE
      port map(D => \InternalDataFromMem\(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(6));
    
    memoryrff_136 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_136, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_136);
    
    memorya49 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya37_2_Z, B => InternalAddr2Memory(8), C
         => memorya51_6_Z, D => memorya369_1_Z, Y => memorya49_Z);
    
    memorya209 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya369_1_Z, 
        C => memorya336_6_Z, D => memorya482_2_Z, Y => 
        memorya209_Z);
    
    memoryrff_45 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_45, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_45);
    
    memoryrff_447 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_447, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_447);
    
    memorya391 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya379_1_Z, 
        C => memorya391_2_Z, D => memorya391_6_Z, Y => 
        memorya391_Z);
    
    memoryrff_298_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya305_2_Z, B => WriteEnable, C => 
        memorya298_6_Z, D => memorya266_0_Z, Y => memorywre_298);
    
    memoryrff_440_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya440_Z, B => WriteEnable, Y => 
        memorywre_440);
    
    memoryrff_47 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_47, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_47);
    
    memoryrff_390_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya390_Z, B => WriteEnable, Y => 
        memorywre_390);
    
    memory_memory_0_0_sr_RNO_139 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_505, B => memoryro_249, C => 
        memorya505_Z, D => memorya249_Z, Y => memoryror_253);
    
    memoryrff_142_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya142_Z, B => WriteEnable, Y => 
        memorywre_142);
    
    memory_memory_0_0_sr_RNO_130 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_323, B => memoryro_195, C => 
        memorya323_Z, D => memorya195_Z, Y => memoryror_200);
    
    memoryrff_255 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_255, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_255);
    
    memoryrff_398 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_398, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_398);
    
    memorya406 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya102_1_Z, B => InternalAddr2Memory(6), 
        C => memorya342_6_Z, D => memorya403_2_Z, Y => 
        memorya406_Z);
    
    memorya320 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_2_Z, B => InternalAddr2Memory(7), C
         => memorya320_6_Z, D => memorya368_2_Z, Y => 
        memorya320_Z);
    
    memorya174 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya162_2_Z, B => memorya110_5_Z, C => 
        InternalAddr2Memory(8), D => memorya289_4_Z, Y => 
        memorya174_Z);
    
    memoryrff_275 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_275, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_275);
    
    memoryrff_163 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_163, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_163);
    
    memorya304_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya304_4_Z, B => memorya57_3_Z, Y => 
        memorya304_6_Z);
    
    memoryrff_76_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya76_Z, B => WriteEnable, Y => 
        memorywre_76);
    
    memorya458 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya362_1_Z, B => InternalAddr2Memory(5), 
        C => memorya362_6_Z, D => memorya482_2_Z, Y => 
        memorya458_Z);
    
    memorya354 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya354_1_Z, 
        C => memorya354_6_Z, D => memorya368_2_Z, Y => 
        memorya354_Z);
    
    memorya291 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya305_2_Z, B => memorya289_6_Z, C => 
        InternalAddr2Memory(7), D => memorya379_1_Z, Y => 
        memorya291_Z);
    
    memoryrff_399_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya399_Z, B => WriteEnable, Y => 
        memorywre_399);
    
    memorya448 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya353_6_Z, 
        C => memorya370_3_Z, D => memorya482_2_Z, Y => 
        memorya448_Z);
    
    memorya344 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya280_0_Z, B => memorya344_6_Z, C => 
        memorya368_2_Z, Y => memorya344_Z);
    
    memoryrff_142 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_142, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_142);
    
    memoryrff_157_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya157_Z, B => WriteEnable, Y => 
        memorywre_157);
    
    memorya266 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya370_3_Z, B => memorya264_6_Z, C => 
        memorya266_0_Z, Y => memorya266_Z);
    
    memoryrff_137_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya193_2_Z, B => WriteEnable, C => 
        memorya264_6_Z, D => memorya9_0_Z, Y => memorywre_137);
    
    memorya236 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya236_0_Z, B => memorya364_1_Z, C => 
        memorya162_2_Z, D => memorya116_2_Z, Y => memorya236_Z);
    
    memorya428_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya434_2_Z, B => memorya364_1_Z, Y => 
        memorya428_5_Z);
    
    memorya155 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya273_4_Z, 
        C => memorya211_3_Z, D => memorya315_5_Z, Y => 
        memorya155_Z);
    
    \memory_memory_0_0_OLDA_RNIDPT31[17]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(17), C => 
        memory_memory_0_0_OLDA_Z(17), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(17));
    
    memorya385_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(0), Y => memorya385_1_Z);
    
    memory_memory_0_0_sr_RNO_10 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_418, B => memoryror_417, C => 
        memoryror_419, D => memoryror_416, Y => memoryror_488);
    
    memoryrff_53 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_53, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_53);
    
    memorya214 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya86_2_Z, B => memorya102_1_Z, C => 
        memorya211_0_Z, D => memorya162_2_Z, Y => memorya214_Z);
    
    memorya145 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya193_2_Z, B => memorya273_6_Z, C => 
        InternalAddr2Memory(8), D => memorya369_1_Z, Y => 
        memorya145_Z);
    
    memoryrff_337 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_337, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_337);
    
    \memory_memory_0_0_OLDA[12]\ : SLE
      port map(D => \InternalDataFromMem\(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(12));
    
    memoryrff_498 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_498, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_498);
    
    memoryrff_259_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya259_Z, B => WriteEnable, Y => 
        memorywre_259);
    
    memoryrff_239_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya239_Z, B => WriteEnable, Y => 
        memorywre_239);
    
    memoryrff_277_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya277_Z, B => WriteEnable, Y => 
        memorywre_277);
    
    memorya184 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya68_2_Z, C
         => memorya312_4_Z, D => memorya440_5_Z, Y => 
        memorya184_Z);
    
    memoryrff_490_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya490_Z, B => WriteEnable, Y => 
        memorywre_490);
    
    memoryrff_24 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_24, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_24);
    
    memorya474 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya86_2_Z, B => memorya498_6_Z, C => 
        InternalAddr2Memory(5), D => memorya362_1_Z, Y => 
        memorya474_Z);
    
    memorya428 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya364_1_Z, B => InternalAddr2Memory(6), 
        C => memorya364_6_Z, D => memorya434_2_Z, Y => 
        memorya428_Z);
    
    memorya324 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya68_1_Z, C
         => memorya197_6_Z, D => memorya370_3_Z, Y => 
        memorya324_Z);
    
    memoryrff_8_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya57_3_Z, C => 
        memorya8_0_Z, D => memorya4_6_Z, Y => memorywre_8);
    
    memoryrff_29_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya29_Z, B => WriteEnable, Y => 
        memorywre_29);
    
    memoryrff_244 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_244, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_244);
    
    memoryrff_192_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya192_Z, B => WriteEnable, Y => 
        memorywre_192);
    
    memorya102_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(1), B => 
        InternalAddr2Memory(2), Y => memorya102_1_Z);
    
    memory_memory_0_0_sr_RNO_331 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_158, B => memoryro_286, C => 
        memorya286_Z, D => memorya158_Z, Y => memoryror_23);
    
    memoryrff_300 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_300, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_300);
    
    memoryrff_14_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya102_1_Z, C => 
        memorya8_0_Z, D => memorya4_6_Z, Y => memorywre_14);
    
    memorya415 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya415_4_Z, 
        C => memorya403_2_Z, D => memorya463_5_Z, Y => 
        memorya415_Z);
    
    memory_memory_0_0_sr_RNO_121 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_201, B => memoryro_457, C => 
        memorya457_Z, D => memorya201_Z, Y => memoryror_205);
    
    memorya125 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya125_2_Z, B => memorya117_1_Z, C => 
        memorya124_0_Z, D => memorya116_2_Z, Y => memorya125_Z);
    
    memory_memory_0_0_sr_RNO_48 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_182, B => memoryror_183, C => 
        memoryror_180, D => memoryror_181, Y => memoryror_429);
    
    memoryrff_443_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya443_Z, B => WriteEnable, Y => 
        memorywre_443);
    
    memory_memory_0_0_sr_RNO_21 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_208, B => memoryror_211, C => 
        memoryror_210, D => memoryror_209, Y => memoryror_436);
    
    memoryrff_229 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_229, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_229);
    
    memorya306_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya304_4_Z, B => memorya354_3_Z, Y => 
        memorya306_6_Z);
    
    memoryrff_465_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya465_Z, B => WriteEnable, Y => 
        memorywre_465);
    
    memoryrff_173_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya173_Z, B => WriteEnable, Y => 
        memorywre_173);
    
    memoryrff_284_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya284_Z, B => WriteEnable, Y => 
        memorywre_284);
    
    memorya196 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya68_1_Z, C
         => memorya162_2_Z, D => memorya197_6_Z, Y => 
        memorya196_Z);
    
    memoryrff_375_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya375_Z, B => WriteEnable, Y => 
        memorywre_375);
    
    memorya278_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(4), Y => memorya278_2_Z);
    
    memory_memory_0_0_sr_RNO_77 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_35, B => memoryror_34, C => 
        memoryror_33, D => memoryror_32, Y => memoryror_392);
    
    memorya484 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya36_1_Z, B => InternalAddr2Memory(4), C
         => memorya372_6_Z, D => memorya482_2_Z, Y => 
        memorya484_Z);
    
    memoryrff_22_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya102_1_Z, B => WriteEnable, C => 
        memorya20_6_Z, D => memorya16_0_Z, Y => memorywre_22);
    
    memorya505 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(2), B => memorya369_3_Z, 
        C => memorya121_5_Z, D => memorya482_2_Z, Y => 
        memorya505_Z);
    
    memoryrff_59_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya59_Z, B => WriteEnable, Y => 
        memorywre_59);
    
    memorya259 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya379_1_Z, B => InternalAddr2Memory(7), 
        C => memorya257_6_Z, D => memorya379_4_Z, Y => 
        memorya259_Z);
    
    memoryrff_75_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya75_Z, B => WriteEnable, Y => 
        memorywre_75);
    
    memoryrff_126 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_126, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_126);
    
    memorya190 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya318_4_Z, B => InternalAddr2Memory(8), 
        C => memorya126_5_Z, D => memorya434_2_Z, Y => 
        memorya190_Z);
    
    memorya249 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya57_3_Z, C
         => memorya121_5_Z, D => memorya482_2_Z, Y => 
        memorya249_Z);
    
    memoryrff_169 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_169, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_169);
    
    memorya56 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya56_0_Z, B => memorya52_4, C => 
        memorya52_2_Z, D => memorya57_3_Z, Y => memorya56_Z);
    
    memory_memory_0_0_sr_RNO_143 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_509, B => memoryro_141, C => 
        memorya509_Z, D => memorya141_Z, Y => memoryror_246);
    
    memorya53 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya84_3_Z, C
         => memorya52_4, D => memorya373_5_Z, Y => memorya53_Z);
    
    memoryrff_425_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya425_Z, B => WriteEnable, Y => 
        memorywre_425);
    
    memoryrff_133 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_133, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_133);
    
    memoryrff_250_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya250_Z, B => WriteEnable, Y => 
        memorywre_250);
    
    memorya27 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya25_3_Z, C
         => memorya52_4, D => memorya315_5_Z, Y => memorya27_Z);
    
    memoryrff_358 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_358, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_358);
    
    memoryrff_230_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya162_2_Z, C => 
        memorya227_0_Z, D => memorya102_5_Z, Y => memorywre_230);
    
    memorya456 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya77_2_Z, C
         => memorya360_6_Z, D => memorya498_3_Z, Y => 
        memorya456_Z);
    
    memory_memory_0_0_sr_RNO_109 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_234, B => memoryro_378, C => 
        memorya378_Z, D => memorya234_Z, Y => memoryror_236);
    
    memoryrff_378 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_378, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_378);
    
    memorya86 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya68_4_Z, B => memorya86_5_Z, C => 
        InternalAddr2Memory(8), D => memorya102_3_Z, Y => 
        memorya86_Z);
    
    memory_memory_0_0_sr_RNO_100 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_495, B => memoryro_175, C => 
        memorya495_Z, D => memorya175_Z, Y => memoryror_227);
    
    memoryrff_44 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_44, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_44);
    
    memorya446 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya370_3_Z, B => memorya126_5_Z, C => 
        InternalAddr2Memory(6), D => memorya434_2_Z, Y => 
        memorya446_Z);
    
    memorya379 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya116_2_Z, B => memorya315_5_Z, C => 
        InternalAddr2Memory(7), D => memorya379_4_Z, Y => 
        memorya379_Z);
    
    memorya83 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya86_2_Z, B => memorya83_6_Z, C => 
        InternalAddr2Memory(8), D => memorya379_1_Z, Y => 
        memorya83_Z);
    
    memoryrff_402_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya402_Z, B => WriteEnable, Y => 
        memorywre_402);
    
    memoryrff_493_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya493_Z, B => WriteEnable, Y => 
        memorywre_493);
    
    memoryrff_52_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya52_Z, B => WriteEnable, Y => 
        memorywre_52);
    
    memoryrff_212 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_212, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_212);
    
    memoryrff_245 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_245, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_245);
    
    memorya362_1 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(1), Y => memorya362_1_Z);
    
    memory_memory_0_0_sr_RNO_322 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_35, B => memoryro_483, C => 
        memorya483_Z, D => memorya35, Y => memoryror_40);
    
    memory_memory_0_0_sr_RNO_276 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_74, B => memoryro_458, C => 
        memorya458_Z, D => memorya74_Z, Y => memoryror_60);
    
    \memory_memory_0_0_OLDA[15]\ : SLE
      port map(D => \InternalDataFromMem\(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(15));
    
    memoryrff_484_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya484_Z, B => WriteEnable, Y => 
        memorywre_484);
    
    memoryrff_18 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_18, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_18);
    
    memoryrff_52 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_52, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_52);
    
    memoryrff_458 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_458, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_458);
    
    memoryrff_327 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_327, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_327);
    
    memorya28 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya29_3_Z, B => memorya364_1_Z, C => 
        memorya52_4, D => memorya16_0_Z, Y => memorya28_Z);
    
    memorya426 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya362_1_Z, B => InternalAddr2Memory(6), 
        C => memorya362_6_Z, D => memorya434_2_Z, Y => 
        memorya426_Z);
    
    memory_memory_0_0_sr_RNO_75 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_2, B => memoryror_0, C => 
        memoryror_1, D => memoryror_3, Y => memoryror_384);
    
    memoryrff_478 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_478, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_478);
    
    memoryrff_6 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_6, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_6);
    
    memoryrff_253_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya253_Z, B => WriteEnable, Y => 
        memorywre_253);
    
    memoryrff_233_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya233_Z, B => WriteEnable, Y => 
        memorywre_233);
    
    memorya389 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya117_1_Z, 
        C => memorya197_6_Z, D => memorya498_3_Z, Y => 
        memorya389_Z);
    
    memoryrff_385 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_385, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_385);
    
    memorya415_4 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(5), Y => memorya415_4_Z);
    
    memoryrff_469 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_469, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_469);
    
    memoryrff_448_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya448_Z, B => WriteEnable, Y => 
        memorywre_448);
    
    memoryrff_16_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya57_3_Z, B => WriteEnable, C => 
        memorya20_6_Z, D => memorya16_0_Z, Y => memorywre_16);
    
    memory_memory_0_0_sr_RNO_301 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_142, B => memoryro_270, C => 
        memorya270_Z, D => memorya142_Z, Y => memoryror_7);
    
    memoryrff_389 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_389, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_389);
    
    memoryrff_241_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya193_2_Z, B => WriteEnable, C => 
        memorya369_5_Z, D => memorya3_0_Z, Y => memorywre_241);
    
    memory_memory_0_0_sr_RNO_247 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_105, B => memoryro_361, C => 
        memorya361_Z, D => memorya105_Z, Y => memoryror_109);
    
    memorya121_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya54_2_Z, B => memorya121_1_Z, Y => 
        memorya121_5_Z);
    
    memory_memory_0_0_sr_RNO_232 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_326, B => memoryro_70, C => 
        memorya326_Z, D => memorya70_Z, Y => memoryror_74);
    
    memory_memory_0_0_sr_RNO_196 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_205, B => memoryro_429, C => 
        memorya429_Z, D => memorya205_Z, Y => memoryror_182);
    
    memoryrff_91 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_91, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_91);
    
    memoryrff_3 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_3, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_3);
    
    memoryrff_88 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_88, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_88);
    
    memoryrff_299 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_299, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_299);
    
    memorya381_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya117_1_Z, B => memorya125_2_Z, Y => 
        memorya381_5_Z);
    
    memorya471 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya487_4_Z, 
        C => memorya482_2_Z, D => memorya503_5_Z, Y => 
        memorya471_Z);
    
    memorya355_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya379_4_Z, B => memorya68_3_Z, Y => 
        memorya355_6_Z);
    
    memoryrff_343_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya343_Z, B => WriteEnable, Y => 
        memorywre_343);
    
    memorya378 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya354_3_Z, 
        C => memorya368_2_Z, D => memorya378_5_Z, Y => 
        memorya378_Z);
    
    memoryrff_139 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_139, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_139);
    
    memorya35_0 : CFG3
      generic map(INIT => x"04")

      port map(A => InternalAddr2Memory(2), B => 
        InternalAddr2Memory(5), C => InternalAddr2Memory(8), Y
         => memorya35_0_Z);
    
    memorya223_0 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(5), Y => memorya223_0_Z);
    
    memorya338_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya20_3_Z, B => memorya354_3_Z, Y => 
        memorya338_6_Z);
    
    memoryrff_196 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_196, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_196);
    
    memorya348_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya86_2_Z, B => memorya364_1_Z, Y => 
        memorya348_5_Z);
    
    memory_memory_0_0_sr_RNO_256 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_366, B => memoryro_238, C => 
        memorya366_Z, D => memorya238_Z, Y => memoryror_103);
    
    memory_memory_0_0_sr_RNO_166 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_232, B => memoryro_280, C => 
        memorya280_Z, D => memorya232_Z, Y => memoryror_159);
    
    memoryrff_374_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya374_Z, B => WriteEnable, Y => 
        memorywre_374);
    
    memoryrff_123 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_123, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_123);
    
    memoryrff_218 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_218, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_218);
    
    memoryrff_306_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya306_Z, B => WriteEnable, Y => 
        memorywre_306);
    
    memory_memory_0_0_sr_RNO_67 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_122, B => memoryror_123, C => 
        memoryror_121, D => memoryror_120, Y => memoryror_414);
    
    memoryrff_507 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_507, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_507);
    
    memoryrff_498_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya498_Z, B => WriteEnable, Y => 
        memorywre_498);
    
    memorya257_0 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(0), Y => memorya257_0_Z);
    
    memorya97 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya117_3_Z, B => memorya98_6_Z, C => 
        InternalAddr2Memory(8), D => memorya353_1_Z, Y => 
        memorya97_Z);
    
    \memory_memory_0_0_OLDA[14]\ : SLE
      port map(D => \InternalDataFromMem\(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(14));
    
    memorya310 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya304_4_Z, B => InternalAddr2Memory(7), 
        C => memorya118_5_Z, D => memorya370_3_Z, Y => 
        memorya310_Z);
    
    memory_memory_0_0_sr_RNO_198 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_380, B => memoryro_188, C => 
        memorya380_Z, D => memorya188_Z, Y => memoryror_180);
    
    memoryrff_148_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya148_Z, B => WriteEnable, Y => 
        memorywre_148);
    
    memoryrff_10 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_10, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_10);
    
    memorya481 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya368_4_Z, B => InternalAddr2Memory(4), 
        C => memorya481_5_Z, D => memorya369_3_Z, Y => 
        memorya481_Z);
    
    memoryrff_71_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya71_Z, B => WriteEnable, Y => 
        memorywre_71);
    
    memoryrff_502 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_502, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_502);
    
    memoryrff_291_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya291_Z, B => WriteEnable, Y => 
        memorywre_291);
    
    memoryrff_184_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya184_Z, B => WriteEnable, Y => 
        memorywre_184);
    
    memorya388 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya197_6_Z, B => memorya370_3_Z, C => 
        InternalAddr2Memory(6), D => memorya391_2_Z, Y => 
        memorya388_Z);
    
    memorya167 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya167_3_Z, 
        C => memorya289_4_Z, D => memorya487_5_Z, Y => 
        memorya167_Z);
    
    memoryrff_412_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya412_Z, B => WriteEnable, Y => 
        memorywre_412);
    
    memoryrff_348 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_348, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_348);
    
    memoryrff_267_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya267_Z, B => WriteEnable, Y => 
        memorywre_267);
    
    memoryrff_501 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_501, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_501);
    
    memory_memory_0_0_sr_RNO_229 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_187, B => memoryro_315, C => 
        memorya315_Z, D => memorya187_Z, Y => memoryror_69);
    
    memory_memory_0_0_sr_RNO_225 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_351, B => memoryro_95, C => 
        memorya351_Z, D => memorya95_Z, Y => memoryror_83);
    
    \memory_memory_0_0_OLDA[10]\ : SLE
      port map(D => \InternalDataFromMem\(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(10));
    
    memoryrff_393_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya393_Z, B => WriteEnable, Y => 
        memorywre_393);
    
    memoryrff_305 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_305, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_305);
    
    memorya57_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(1), B => 
        InternalAddr2Memory(2), Y => memorya57_3_Z);
    
    memory_memory_0_0_sr_RNO_168 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_107, B => memoryro_411, C => 
        memorya411_Z, D => memorya107_Z, Y => memoryror_149);
    
    memoryrff_15_RNO : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya463_5_Z, B => memorya4_6_Z, C => 
        InternalAddr2Memory(8), D => WriteEnable, Y => 
        memorywre_15);
    
    memorya236_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya45_3_Z, B => InternalAddr2Memory(8), Y
         => memorya236_0_Z);
    
    memoryrff_181_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya181_Z, B => WriteEnable, Y => 
        memorywre_181);
    
    memorya194 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya66_1_Z, C
         => memorya162_2_Z, D => memorya320_6_Z, Y => 
        memorya194_Z);
    
    memoryrff_59 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_59, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_59);
    
    memoryrff_397 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_397, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_397);
    
    memoryrff_309 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_309, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_309);
    
    memoryrff_285_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya285_Z, B => WriteEnable, Y => 
        memorywre_285);
    
    memoryrff_439 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_439, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_439);
    
    memorya98 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya84_2_Z, B => memorya98_6_Z, C => 
        InternalAddr2Memory(8), D => memorya354_1_Z, Y => 
        memorya98_Z);
    
    memoryrff_185_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya185_Z, B => WriteEnable, Y => 
        memorywre_185);
    
    memorya418 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya354_1_Z, 
        C => memorya354_6_Z, D => memorya498_3_Z, Y => 
        memorya418_Z);
    
    memorya314 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya312_4_Z, B => InternalAddr2Memory(7), 
        C => memorya370_3_Z, D => memorya378_5_Z, Y => 
        memorya314_Z);
    
    memoryrff_80 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_80, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_80);
    
    memoryrff_227_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya227_Z, B => WriteEnable, Y => 
        memorywre_227);
    
    memoryrff_163_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya163_Z, B => WriteEnable, Y => 
        memorywre_163);
    
    memoryrff_506_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya506_Z, B => WriteEnable, Y => 
        memorywre_506);
    
    memoryrff_282_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya282_Z, B => WriteEnable, Y => 
        memorywre_282);
    
    memoryrff_448 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_448, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_448);
    
    memoryrff_365_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya365_Z, B => WriteEnable, Y => 
        memorywre_365);
    
    memory_memory_0_0_sr_RNO_97 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_398, B => memoryro_94, C => 
        memorya398_Z, D => memorya94_Z, Y => memoryror_215);
    
    memorya362 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya362_1_Z, 
        C => memorya116_2_Z, D => memorya362_6_Z, Y => 
        memorya362_Z);
    
    memorya332 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya204_6_Z, B => memorya368_2_Z, C => 
        memorya268_0_Z, Y => memorya332_Z);
    
    memorya169 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya121_1_Z, B => InternalAddr2Memory(8), 
        C => memorya296_6_Z, D => memorya434_2_Z, Y => 
        memorya169_Z);
    
    memoryrff_198_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya198_Z, B => WriteEnable, Y => 
        memorywre_198);
    
    memorya278 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya102_1_Z, 
        C => memorya278_2_Z, D => memorya278_6_Z, Y => 
        memorya278_Z);
    
    memory_memory_0_0_sr_RNO_65 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_127, B => memoryror_125, C => 
        memoryror_124, D => memoryror_126, Y => memoryror_415);
    
    memoryrff_446_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya446_Z, B => WriteEnable, Y => 
        memorywre_446);
    
    memorya139 : CFG3
      generic map(INIT => x"20")

      port map(A => memorya264_6_Z, B => InternalAddr2Memory(8), 
        C => memorya395_5_Z, Y => memorya139_Z);
    
    memorya115 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya67_2_Z, C
         => memorya116_4_Z, D => memorya499_5_Z, Y => 
        memorya115_Z);
    
    memoryrff_93_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya93_Z, B => WriteEnable, Y => 
        memorywre_93);
    
    memoryrff_33_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya33_Z, B => WriteEnable, Y => 
        memorywre_33);
    
    memoryrff_117 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_117, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_117);
    
    memorya272 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_2_Z, B => InternalAddr2Memory(7), C
         => memorya273_6_Z, D => memorya278_2_Z, Y => 
        memorya272_Z);
    
    memoryrff_504 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_504, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_504);
    
    memoryrff_259 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_259, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_259);
    
    memoryrff_342_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya342_Z, B => WriteEnable, Y => 
        memorywre_342);
    
    memory_memory_0_0_sr_RNO_234 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_325, B => memoryro_69, C => 
        memorya325_Z, D => memorya69_Z, Y => memoryror_75);
    
    memory_memory_0_0_sr_RNO_19 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_388, B => memoryror_389, C => 
        memoryror_391, D => memoryror_390, Y => memoryror_481);
    
    memorya487_4 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(3), Y => memorya487_4_Z);
    
    memorya494 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(4), B => memorya370_3_Z, 
        C => memorya110_5_Z, D => memorya482_2_Z, Y => 
        memorya494_Z);
    
    memorya469 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya84_3_Z, B => InternalAddr2Memory(5), C
         => memorya213_5_Z, D => memorya498_3_Z, Y => 
        memorya469_Z);
    
    memorya363 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya41_3_Z, B => InternalAddr2Memory(7), C
         => memorya299_5_Z, D => memorya368_2_Z, Y => 
        memorya363_Z);
    
    memoryrff_279 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_279, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_279);
    
    memory_memory_0_0_sr_RNO_37 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_161, B => memoryror_163, C => 
        memoryror_162, D => memoryror_160, Y => memoryror_424);
    
    memory_memory_0_0_sr_RNO_172 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_389, B => memoryro_165, C => 
        memorya389_Z, D => memorya165_Z, Y => memoryror_155);
    
    memoryrff_28_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya28_Z, B => WriteEnable, Y => 
        memorywre_28);
    
    memoryrff_123_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya121_4_Z, C => 
        memorya315_5_Z, D => memorya111_0_Z, Y => memorywre_123);
    
    memorya439 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya487_4_Z, 
        C => memorya434_2_Z, D => memorya503_5_Z, Y => 
        memorya439_Z);
    
    memorya333 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya77_2_Z, B => memorya333_6_Z, C => 
        InternalAddr2Memory(7), D => memorya117_1_Z, Y => 
        memorya333_Z);
    
    memory_memory_0_0_sr_RNO_54 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_87, B => memoryror_84, C => 
        memoryror_86, D => memoryror_85, Y => memoryror_405);
    
    memory_memory_0_0_sr_RNO_202 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_137, B => memoryro_425, C => 
        memorya425_Z, D => memorya137, Y => memoryror_189);
    
    memoryrff_313 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_313, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_313);
    
    memoryrff_129 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_129, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_129);
    
    memoryrff_325_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya325_Z, B => WriteEnable, Y => 
        memorywre_325);
    
    memory_memory_0_0_sr_RNO_135 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_511, B => memoryro_191, C => 
        memorya511_Z, D => memorya191_Z, Y => memoryror_243);
    
    memoryrff_156 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_156, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_156);
    
    memorya98_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya102_4_Z, B => memorya368_4_Z, Y => 
        memorya98_6_Z);
    
    memoryrff_177_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya177_Z, B => WriteEnable, Y => 
        memorywre_177);
    
    memory_memory_0_0_sr_RNO_335 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_106, B => memoryro_490, C => 
        memorya490_Z, D => memorya106_Z, Y => memoryror_28);
    
    memoryrff_27_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya27_Z, B => WriteEnable, Y => 
        memorywre_27);
    
    memory_memory_0_0_sr_RNO_231 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_44, B => memoryro_460, C => 
        memorya460_Z, D => memorya44, Y => memoryror_68);
    
    memory_memory_0_0_sr_RNO_16 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_399, B => memoryror_396, C => 
        memoryror_397, D => memoryror_398, Y => memoryror_483);
    
    memoryrff_176 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_176, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_176);
    
    memorya68_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(5), Y => memorya68_4_Z);
    
    memorya288 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_2_Z, B => InternalAddr2Memory(7), C
         => memorya289_6_Z, D => memorya305_2_Z, Y => 
        memorya288_Z);
    
    memoryrff_193 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_193, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_193);
    
    memory_memory_0_0_sr_RNO_230 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_77, B => memoryro_333, C => 
        memorya333_Z, D => memorya77_Z, Y => memoryror_70);
    
    memory_memory_0_0_sr_RNO_84 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_471, B => memoryro_135, C => 
        memorya471_Z, D => memorya135_Z, Y => memoryror_222);
    
    memorya282 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya354_3_Z, B => memorya273_4_Z, C => 
        memorya278_2_Z, D => memorya266_0_Z, Y => memorya282_Z);
    
    memory_memory_0_0_sr_RNO_343 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya3_0_Z, B => memorya369_5_Z, C => 
        memorya193_2_Z, Y => memorya241);
    
    memoryrff_316_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya316_Z, B => WriteEnable, Y => 
        memorywre_316);
    
    memoryrff_279_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya279_Z, B => WriteEnable, Y => 
        memorywre_279);
    
    memorya336_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya20_3_Z, B => memorya57_3_Z, Y => 
        memorya336_6_Z);
    
    memorya29_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(1), Y => memorya29_3_Z);
    
    memoryrff_69_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya69_Z, B => WriteEnable, Y => 
        memorywre_69);
    
    memoryrff_58_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya58_Z, B => WriteEnable, Y => 
        memorywre_58);
    
    memoryrff_496_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya496_Z, B => WriteEnable, Y => 
        memorywre_496);
    
    memory_memory_0_0_sr_RNO_95 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_214, B => memoryro_390, C => 
        memorya390_Z, D => memorya214_Z, Y => memoryror_218);
    
    memorya118_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya54_2_Z, B => memorya102_1_Z, Y => 
        memorya118_5_Z);
    
    memorya45_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya52_4, B => memorya45_3_Z, Y => 
        memorya45_6_Z);
    
    memorya219 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya25_3_Z, B => InternalAddr2Memory(8), C
         => memorya315_5_Z, D => memorya482_2_Z, Y => 
        memorya219_Z);
    
    memoryrff_392_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya392_Z, B => WriteEnable, Y => 
        memorywre_392);
    
    memoryrff_280 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_280, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_280);
    
    memory_memory_0_0_sr_RNO_71 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_58, B => memoryror_59, C => 
        memoryror_57, D => memoryror_56, Y => memoryror_398);
    
    memory_memory_0_0_sr_RNO_5 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_440, B => memoryror_441, C => 
        memoryror_443, D => memoryror_442, Y => memoryror_494);
    
    memoryrff_57_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya57_Z, B => WriteEnable, Y => 
        memorywre_57);
    
    memoryrff_208_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya208_Z, B => WriteEnable, Y => 
        memorywre_208);
    
    memorya29 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya29_3_Z, C
         => memorya52_4, D => memorya381_5_Z, Y => memorya29_Z);
    
    memoryrff_300_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya300_Z, B => WriteEnable, Y => 
        memorywre_300);
    
    memoryrff_55 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_55, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_55);
    
    memorya121_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(2), Y => memorya121_4_Z);
    
    memory_memory_0_0_sr_RNO_35 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_248, B => memoryror_249, C => 
        memoryror_251, D => memoryror_250, Y => memoryror_446);
    
    memory_memory_0_0_sr_RNO_152 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_161, B => memoryro_289, C => 
        memorya289_Z, D => memorya161_Z, Y => memoryror_161);
    
    memoryrff_357 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_357, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_357);
    
    memorya399 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya4_3_Z, B => InternalAddr2Memory(6), C
         => memorya463_5_Z, D => memorya498_3_Z, Y => 
        memorya399_Z);
    
    memory_memory_0_0_sr_RNO_123 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_346, B => memoryro_202, C => 
        memorya346_Z, D => memorya202_Z, Y => memoryror_204);
    
    memoryrff_341_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya341_Z, B => WriteEnable, Y => 
        memorywre_341);
    
    memorya416 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya353_6_Z, B => memorya370_3_Z, C => 
        InternalAddr2Memory(6), D => memorya434_2_Z, Y => 
        memorya416_Z);
    
    memoryrff_57 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_57, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_57);
    
    memoryrff_429 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_429, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_429);
    
    memoryrff_377 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_377, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_377);
    
    memory_memory_0_0_sr_RNO_199 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_427, B => memoryro_75, C => 
        memorya427_Z, D => memorya75_Z, Y => memoryror_181);
    
    memoryrff_76 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_76, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_76);
    
    memory_memory_0_0_sr_RNO_190 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_391, B => memoryro_215, C => 
        memorya391_Z, D => memorya215_Z, Y => memoryror_142);
    
    memoryrff_62_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya62_Z, B => WriteEnable, Y => 
        memorywre_62);
    
    memory_memory_0_0_sr_RNO_278 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_72, B => memoryro_504, C => 
        memorya504_Z, D => memorya72_Z, Y => memoryror_63);
    
    memory_memory_0_0_sr_RNO_8 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_426, B => memoryror_424, C => 
        memoryror_427, D => memoryror_425, Y => memoryror_490);
    
    memoryrff_482 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_482, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_482);
    
    memoryrff_309_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya309_Z, B => WriteEnable, Y => 
        memorywre_309);
    
    memoryrff_484 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_484, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_484);
    
    memory_memory_0_0_sr_RNO_137 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_250, B => memoryro_362, C => 
        memorya362_Z, D => memorya250_Z, Y => memoryror_252);
    
    memoryrff_263 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_263, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_263);
    
    memoryrff_11_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya11_Z, B => WriteEnable, Y => 
        memorywre_11);
    
    \memory_memory_0_0_OLDA_RNI7KU31[20]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(20), C => 
        memory_memory_0_0_OLDA_Z(20), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(20));
    
    memoryrff_311 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_311, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_311);
    
    memorya400 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya336_6_Z, B => memorya370_3_Z, C => 
        InternalAddr2Memory(6), D => memorya403_2_Z, Y => 
        memorya400_Z);
    
    memoryrff_286_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya286_Z, B => WriteEnable, Y => 
        memorywre_286);
    
    memory_memory_0_0_sr_RNO_169 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_30, B => memoryro_494, C => 
        memorya494_Z, D => memorya30_Z, Y => memoryror_151);
    
    memoryrff_270_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya270_Z, B => WriteEnable, Y => 
        memorywre_270);
    
    memory_memory_0_0_sr_RNO_160 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_46, B => memoryro_478, C => 
        memorya478_Z, D => memorya46_Z, Y => memoryror_167);
    
    memoryrff_115 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_115, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_115);
    
    memorya3_0 : CFG2
      generic map(INIT => x"2")

      port map(A => memorya368_4_Z, B => InternalAddr2Memory(8), 
        Y => memorya3_0_Z);
    
    memory_memory_0_0_sr_RNO_216 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_341, B => memoryro_85, C => 
        memorya341_Z, D => memorya85_Z, Y => memoryror_91);
    
    memoryrff_94_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya94_Z, B => WriteEnable, Y => 
        memorywre_94);
    
    memoryrff_364_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya364_Z, B => WriteEnable, Y => 
        memorywre_364);
    
    memoryrff_34_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya354_1_Z, B => WriteEnable, C => 
        memorya36_6_Z, D => memorya10_0_Z, Y => memorywre_34);
    
    memoryrff_382 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_382, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_382);
    
    memorya305_2 : CFG2
      generic map(INIT => x"8")

      port map(A => InternalAddr2Memory(8), B => 
        InternalAddr2Memory(5), Y => memorya305_2_Z);
    
    memory_memory_0_0_sr_RNO_204 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_338, B => memoryro_50, C => 
        memorya338_Z, D => memorya50_Z, Y => memoryror_176);
    
    memoryrff_400_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya400_Z, B => WriteEnable, Y => 
        memorywre_400);
    
    memory_memory_0_0_sr_RNO_186 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_14, B => memoryro_510, C => 
        memorya510_Z, D => memorya14, Y => memoryror_135);
    
    memoryrff_199 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_199, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_199);
    
    memoryrff_102_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya102_Z, B => WriteEnable, Y => 
        memorywre_102);
    
    \memory_memory_0_0_OLDA[4]\ : SLE
      port map(D => \InternalDataFromMem\(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(4));
    
    memoryrff_249 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_249, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_249);
    
    memoryrff_391_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya391_Z, B => WriteEnable, Y => 
        memorywre_391);
    
    memory_memory_0_0_sr_RNO_105 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_507, B => memoryro_59, C => 
        memorya507_Z, D => memorya59_Z, Y => memoryror_229);
    
    memory_memory_0_0_sr_RNO_377 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya36_6_Z, B => memorya379_1_Z, C => 
        memorya35_0_Z, Y => memorya35);
    
    memoryrff_386 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_386, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_386);
    
    memorya102_3 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(3), B => 
        InternalAddr2Memory(0), Y => memorya102_3_Z);
    
    memory_memory_0_0_sr_RNO_305 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_130, B => memoryro_450, C => 
        memorya450_Z, D => memorya130_Z, Y => memoryror_0);
    
    memoryrff_153 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_153, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_153);
    
    memory_memory_0_0_sr_RNO_201 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_231, B => memoryro_439, C => 
        memorya439_Z, D => memorya231_Z, Y => memoryror_190);
    
    memoryrff_200 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_200, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_200);
    
    \memory_memory_0_0_OLDA[23]\ : SLE
      port map(D => \InternalDataFromMem\(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(23));
    
    memory_memory_0_0_sr_RNO_340 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya83_6_Z, B => memorya86_2_Z, C => 
        memorya20_0_Z, Y => memorya80);
    
    memoryrff_324_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya324_Z, B => WriteEnable, Y => 
        memorywre_324);
    
    memorya491 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(4), B => memorya379_4_Z, 
        C => memorya299_5_Z, D => memorya482_2_Z, Y => 
        memorya491_Z);
    
    memorya304_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(3), Y => memorya304_4_Z);
    
    memoryrff_173 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_173, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_173);
    
    memoryrff_146 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_146, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_146);
    
    memory_memory_0_0_sr_RNO_273 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_117, B => memoryro_373, C => 
        memorya373_Z, D => memorya117_Z, Y => memoryror_123);
    
    memory_memory_0_0_sr_RNO_258 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_12, B => memoryro_492, C => 
        memorya492_Z, D => memorya12, Y => memoryror_100);
    
    memoryrff_487 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_487, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_487);
    
    memorya398 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya4_3_Z, B => InternalAddr2Memory(6), C
         => memorya142_5_Z, D => memorya370_3_Z, Y => 
        memorya398_Z);
    
    memorya36_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya52_4, B => memorya68_3_Z, Y => 
        memorya36_6_Z);
    
    memory_memory_0_0_sr_RNO_227 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_210, B => memoryro_434, C => 
        memorya434_Z, D => memorya210_Z, Y => memoryror_80);
    
    memory_memory_0_0_sr_RNO_200 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_312, B => memoryro_200, C => 
        memorya312_Z, D => memorya200_Z, Y => memoryror_191);
    
    memoryrff_273_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya273_Z, B => WriteEnable, Y => 
        memorywre_273);
    
    memorya37 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya37_2_Z, B => InternalAddr2Memory(8), C
         => memorya36_6_Z, D => memorya117_1_Z, Y => memorya37_Z);
    
    memory_memory_0_0_sr_RNO_361 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya45_6_Z, B => memorya52_2_Z, C => 
        memorya12_0_Z, Y => memorya44);
    
    memorya365 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya45_3_Z, B => InternalAddr2Memory(7), C
         => memorya45_5_Z, D => memorya368_2_Z, Y => memorya365_Z);
    
    \memory_memory_0_0_OLDA[30]\ : SLE
      port map(D => \InternalDataFromMem\(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memory_memory_0_0_OLDA_Z(30));
    
    memorya335 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya4_3_Z, C
         => memorya368_2_Z, D => memorya463_5_Z, Y => 
        memorya335_Z);
    
    memory_memory_0_0_sr_RNO_188 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_314, B => memoryro_138, C => 
        memorya314_Z, D => memorya138, Y => memoryror_140);
    
    memoryrff_452_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya452_Z, B => WriteEnable, Y => 
        memorywre_452);
    
    memoryrff_413 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_413, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_413);
    
    memoryrff_410 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_410, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_410);
    
    memoryrff_432_RNO : CFG3
      generic map(INIT => x"80")

      port map(A => memorya432_0_Z, B => WriteEnable, C => 
        memorya368_6_Z, Y => memorywre_432);
    
    memoryrff_402 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_402, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_402);
    
    memorya197_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya4_3_Z, B => memorya84_3_Z, Y => 
        memorya197_6_Z);
    
    memoryrff_218_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya218_Z, B => WriteEnable, Y => 
        memorywre_218);
    
    memoryrff_61 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_61, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_61);
    
    memoryrff_73 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_73, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_73);
    
    memoryrff_404 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_404, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_404);
    
    memorya99 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya116_2_Z, B => memorya98_6_Z, C => 
        InternalAddr2Memory(8), D => memorya379_1_Z, Y => 
        memorya99_Z);
    
    memoryrff_310_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya310_Z, B => WriteEnable, Y => 
        memorywre_310);
    
    memoryrff_182 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_182, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_182);
    
    memoryrff_186_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya186_Z, B => WriteEnable, Y => 
        memorywre_186);
    
    memoryrff_114 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_114, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_114);
    
    \memory_memory_0_0_OLDA_RNIFSU31[28]\ : CFG4
      generic map(INIT => x"50D8")

      port map(A => memory_memory_0_0_en_Z, B => 
        memory_memory_0_0_NEWA(28), C => 
        memory_memory_0_0_OLDA_Z(28), D => memory_memory_0_0_sr_Z, 
        Y => \InternalDataFromMem\(28));
    
    memory_memory_0_0_sr_RNO_61 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_106, B => memoryror_105, C => 
        memoryror_104, D => memoryror_107, Y => memoryror_410);
    
    memory_memory_0_0_sr_RNO_131 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_469, B => memoryro_229, C => 
        memorya469_Z, D => memorya229, Y => memoryror_203);
    
    memoryrff_499 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_499, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_499);
    
    memoryrff_233 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_233, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_233);
    
    memorya378_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya54_2_Z, B => memorya362_1_Z, Y => 
        memorya378_5_Z);
    
    memoryrff_403_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya403_Z, B => WriteEnable, Y => 
        memorywre_403);
    
    memorya38 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya52_2_Z, B => InternalAddr2Memory(8), C
         => memorya36_6_Z, D => memorya102_1_Z, Y => memorya38_Z);
    
    memoryrff_54 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_54, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_54);
    
    memoryrff_319_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya319_Z, B => WriteEnable, Y => 
        memorywre_319);
    
    memoryrff_302 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_302, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_302);
    
    memory_memory_0_0_sr_RNO_357 : CFG3
      generic map(INIT => x"20")

      port map(A => memorya4_6_Z, B => InternalAddr2Memory(8), C
         => memorya368_6_Z, Y => memorya0);
    
    memoryrff_347 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_347, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_347);
    
    memoryrff_244_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya244_Z, B => WriteEnable, Y => 
        memorywre_244);
    
    memorya13 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya13_0_Z, B => InternalAddr2Memory(8), C
         => memorya117_1_Z, D => memorya4_6_Z, Y => memorya13_Z);
    
    memorya102_4 : CFG2
      generic map(INIT => x"1")

      port map(A => InternalAddr2Memory(7), B => 
        InternalAddr2Memory(4), Y => memorya102_4_Z);
    
    memorya345_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya369_3_Z, B => memorya25_3_Z, Y => 
        memorya345_6_Z);
    
    memoryrff_31 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_31, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_31);
    
    memorya450 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya66_1_Z, C
         => memorya354_6_Z, D => memorya498_3_Z, Y => 
        memorya450_Z);
    
    memoryrff_28 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_28, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_28);
    
    memorya440_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya434_2_Z, B => memorya125_2_Z, Y => 
        memorya440_5_Z);
    
    memorya440 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya125_2_Z, B => InternalAddr2Memory(6), 
        C => memorya376_6_Z, D => memorya434_2_Z, Y => 
        memorya440_Z);
    
    memory_memory_0_0_sr_RNO_253 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_386, B => memoryro_226, C => 
        memorya386_Z, D => memorya226_Z, Y => memoryror_96);
    
    memory_memory_0_0_sr_RNO_107 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_110, B => memoryro_430, C => 
        memorya430_Z, D => memorya110_Z, Y => memoryror_231);
    
    memoryrff_284 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_284, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_284);
    
    memoryrff_167_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya167_Z, B => WriteEnable, Y => 
        memorywre_167);
    
    memorya472 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(5), B => memorya125_2_Z, 
        C => memorya376_6_Z, D => memorya482_2_Z, Y => 
        memorya472_Z);
    
    memoryrff_306 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_306, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_306);
    
    memorya37_2 : CFG2
      generic map(INIT => x"2")

      port map(A => InternalAddr2Memory(5), B => 
        InternalAddr2Memory(1), Y => memorya37_2_Z);
    
    memory_memory_0_0_sr_RNO_348 : CFG3
      generic map(INIT => x"80")

      port map(A => memorya503_5_Z, B => memorya111_0_Z, C => 
        memorya167_3_Z, Y => memorya247);
    
    memoryrff_96_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya96_Z, B => WriteEnable, Y => 
        memorywre_96);
    
    memoryrff_36_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya36_1_Z, B => WriteEnable, C => 
        memorya36_6_Z, D => memorya20_0_Z, Y => memorywre_36);
    
    memoryrff_159 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_159, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_159);
    
    memorya260 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya68_2_Z, B => InternalAddr2Memory(7), C
         => memorya257_6_Z, D => memorya260_1_Z, Y => 
        memorya260_Z);
    
    memoryrff_410_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya410_Z, B => WriteEnable, Y => 
        memorywre_410);
    
    memoryrff_407 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_407, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_407);
    
    memoryrff_269_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya264_1_Z, B => WriteEnable, C => 
        memorya268_6_Z, D => memorya261_0_Z, Y => memorywre_269);
    
    memory_memory_0_0_sr_RNO_18 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_393, B => memoryror_392, C => 
        memoryror_395, D => memoryror_394, Y => memoryror_482);
    
    memoryrff_179 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_179, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_179);
    
    memorya124_0 : CFG3
      generic map(INIT => x"01")

      port map(A => InternalAddr2Memory(1), B => 
        InternalAddr2Memory(7), C => InternalAddr2Memory(8), Y
         => memorya124_0_Z);
    
    memoryrff_112_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya112_Z, B => WriteEnable, Y => 
        memorywre_112);
    
    memorya376 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(7), B => memorya125_2_Z, 
        C => memorya116_2_Z, D => memorya376_6_Z, Y => 
        memorya376_Z);
    
    memoryrff_216 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_216, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_216);
    
    memoryrff_127_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya127_Z, B => WriteEnable, Y => 
        memorywre_127);
    
    memorya77 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(8), B => memorya45_3_Z, C
         => memorya68_4_Z, D => memorya77_5_Z, Y => memorya77_Z);
    
    memorya420 : CFG4
      generic map(INIT => x"4000")

      port map(A => InternalAddr2Memory(6), B => memorya36_1_Z, C
         => memorya356_6_Z, D => memorya498_3_Z, Y => 
        memorya420_Z);
    
    memorya292 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya36_1_Z, B => InternalAddr2Memory(7), C
         => memorya292_6_Z, D => memorya370_3_Z, Y => 
        memorya292_Z);
    
    memory_memory_0_0_sr_RNO_91 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_337, B => memoryro_209, C => 
        memorya337_Z, D => memorya209_Z, Y => memoryror_209);
    
    memoryrff_481_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya481_Z, B => WriteEnable, Y => 
        memorywre_481);
    
    memorya4_6 : CFG3
      generic map(INIT => x"10")

      port map(A => InternalAddr2Memory(6), B => 
        InternalAddr2Memory(7), C => memorya4_3_Z, Y => 
        memorya4_6_Z);
    
    memorya339_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya379_4_Z, B => memorya20_3_Z, Y => 
        memorya339_6_Z);
    
    memorya482 : CFG4
      generic map(INIT => x"2000")

      port map(A => memorya354_1_Z, B => InternalAddr2Memory(4), 
        C => memorya370_6_Z, D => memorya482_2_Z, Y => 
        memorya482_Z);
    
    memorya299_5 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya379_1_Z, B => memorya45_2_Z, Y => 
        memorya299_5_Z);
    
    memoryrff_294_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya294_Z, B => WriteEnable, Y => 
        memorywre_294);
    
    memorya275 : CFG4
      generic map(INIT => x"0800")

      port map(A => memorya278_2_Z, B => memorya273_6_Z, C => 
        InternalAddr2Memory(7), D => memorya379_1_Z, Y => 
        memorya275_Z);
    
    memoryrff_356_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya356_Z, B => WriteEnable, Y => 
        memorywre_356);
    
    memoryrff_336_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya336_Z, B => WriteEnable, Y => 
        memorywre_336);
    
    memorya68_6 : CFG2
      generic map(INIT => x"8")

      port map(A => memorya68_4_Z, B => memorya68_3_Z, Y => 
        memorya68_6_Z);
    
    memoryrff_229_RNO : CFG4
      generic map(INIT => x"8000")

      port map(A => WriteEnable, B => memorya193_2_Z, C => 
        memorya227_0_Z, D => memorya101_5_Z, Y => memorywre_229);
    
    memory_memory_0_0_sr_RNO_292 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_279, B => memoryro_7, C => 
        memorya279_Z, D => memorya7_Z, Y => memoryror_14);
    
    memoryrff_102 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_102, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_102);
    
    memorya108 : CFG4
      generic map(INIT => x"8000")

      port map(A => memorya364_1_Z, B => memorya102_4_Z, C => 
        memorya116_2_Z, D => memorya20_0_Z, Y => memorya108_Z);
    
    memory_memory_0_0_sr_RNO_332 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => memoryro_472, B => memoryro_104, C => 
        memorya472_Z, D => memorya104_Z, Y => memoryror_31);
    
    memoryrff_444_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya444_Z, B => WriteEnable, Y => 
        memorywre_444);
    
    memoryrff_143 : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        memorywre_143, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => memoryro_143);
    
    memory_memory_0_0_sr_RNO_31 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => memoryror_202, B => memoryror_201, C => 
        memoryror_200, D => memoryror_203, Y => memoryror_434);
    
    memory_memory_0_0_sr_RNO_112 : CFG4
      generic map(INIT => x"EAC0")

      port map(A => memoryro_228, B => memoryro_292, C => 
        memorya292_Z, D => memorya228_Z, Y => memoryror_233);
    
    memoryrff_70_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => memorya70_Z, B => WriteEnable, Y => 
        memorywre_70);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Timestamp is

    port( TimeStampValue     : out   std_logic_vector(31 downto 0);
          getTime            : in    std_logic;
          enableTimestampGen : in    std_logic;
          sb_sb_0_FIC_0_CLK  : in    std_logic;
          resetn_arst        : in    std_logic
        );

end Timestamp;

architecture DEF_ARCH of Timestamp is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal counter_Z : std_logic_vector(31 downto 0);
    signal counter_s : std_logic_vector(30 downto 0);
    signal prescaler_Z : std_logic_vector(5 downto 0);
    signal prescaler_5_Z : std_logic_vector(4 downto 3);
    signal state_Z : std_logic_vector(0 to 0);
    signal counter_s_Z : std_logic_vector(31 to 31);
    signal counter_cry_Z : std_logic_vector(30 downto 1);
    signal counter_cry_Y : std_logic_vector(30 downto 1);
    signal counter_s_FCO : std_logic_vector(31 to 31);
    signal counter_s_Y : std_logic_vector(31 to 31);
    signal \VCC\, un1_prescaler_axbxc0_Z, \GND\, 
        un1_prescaler_axbxc1_Z, un1_prescaler_axbxc2_Z, 
        un1_prescaler_axbxc5_Z, prescaler_2_sqmuxa_Z, 
        state_0_sqmuxa_Z, countere, counter_s_830_FCO, 
        counter_s_830_S, counter_s_830_Y, un1_prescaler_c2, 
        counter_0_sqmuxa_0_Z, un6_enable_3_Z, un1_prescaler_c4
         : std_logic;

begin 


    \timestamp[20]\ : SLE
      port map(D => counter_Z(20), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(20));
    
    \prescaler_5[3]\ : CFG4
      generic map(INIT => x"1230")

      port map(A => un1_prescaler_c2, B => countere, C => 
        prescaler_Z(3), D => prescaler_Z(2), Y => 
        prescaler_5_Z(3));
    
    un1_prescaler_axbxc1 : CFG3
      generic map(INIT => x"6A")

      port map(A => prescaler_Z(1), B => prescaler_Z(0), C => 
        counter_0_sqmuxa_0_Z, Y => un1_prescaler_axbxc1_Z);
    
    \counter_cry[21]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(21), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(20), S => counter_s(21), Y
         => counter_cry_Y(21), FCO => counter_cry_Z(21));
    
    \timestamp[16]\ : SLE
      port map(D => counter_Z(16), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(16));
    
    \counter_cry[18]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(18), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(17), S => counter_s(18), Y
         => counter_cry_Y(18), FCO => counter_cry_Z(18));
    
    \timestamp[22]\ : SLE
      port map(D => counter_Z(22), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(22));
    
    \prescaler[0]\ : SLE
      port map(D => un1_prescaler_axbxc0_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        prescaler_Z(0));
    
    \counter_cry[22]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(22), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(21), S => counter_s(22), Y
         => counter_cry_Y(22), FCO => counter_cry_Z(22));
    
    \counter[24]\ : SLE
      port map(D => counter_s(24), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(24));
    
    \counter[17]\ : SLE
      port map(D => counter_s(17), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(17));
    
    \timestamp[4]\ : SLE
      port map(D => counter_Z(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(4));
    
    \counter[2]\ : SLE
      port map(D => counter_s(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(2));
    
    \counter[7]\ : SLE
      port map(D => counter_s(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(7));
    
    \counter_cry[15]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(15), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(14), S => counter_s(15), Y
         => counter_cry_Y(15), FCO => counter_cry_Z(15));
    
    \counter_s[31]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(31), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(30), S => counter_s_Z(31), Y
         => counter_s_Y(31), FCO => counter_s_FCO(31));
    
    \counter_cry[26]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(26), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(25), S => counter_s(26), Y
         => counter_cry_Y(26), FCO => counter_cry_Z(26));
    
    \timestamp[13]\ : SLE
      port map(D => counter_Z(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(13));
    
    \counter_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => counter_Z(0), Y => counter_s(0));
    
    \counter_cry[20]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(20), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(19), S => counter_s(20), Y
         => counter_cry_Y(20), FCO => counter_cry_Z(20));
    
    \counter[6]\ : SLE
      port map(D => counter_s(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(6));
    
    \timestamp[11]\ : SLE
      port map(D => counter_Z(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(11));
    
    \counter_cry[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(13), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(12), S => counter_s(13), Y
         => counter_cry_Y(13), FCO => counter_cry_Z(13));
    
    \prescaler[5]\ : SLE
      port map(D => un1_prescaler_axbxc5_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        prescaler_Z(5));
    
    \timestamp[24]\ : SLE
      port map(D => counter_Z(24), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(24));
    
    \counter_cry[27]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(27), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(26), S => counter_s(27), Y
         => counter_cry_Y(27), FCO => counter_cry_Z(27));
    
    \timestamp[19]\ : SLE
      port map(D => counter_Z(19), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(19));
    
    \counter[8]\ : SLE
      port map(D => counter_s(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(8));
    
    \counter[22]\ : SLE
      port map(D => counter_s(22), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(22));
    
    un1_prescaler_ac0_5 : CFG3
      generic map(INIT => x"80")

      port map(A => prescaler_Z(2), B => un1_prescaler_c2, C => 
        prescaler_Z(3), Y => un1_prescaler_c4);
    
    \counter[16]\ : SLE
      port map(D => counter_s(16), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(16));
    
    \timestamp[7]\ : SLE
      port map(D => counter_Z(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(7));
    
    un1_prescaler_axbxc2 : CFG2
      generic map(INIT => x"6")

      port map(A => un1_prescaler_c2, B => prescaler_Z(2), Y => 
        un1_prescaler_axbxc2_Z);
    
    \counter_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(6), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(5), S => counter_s(6), Y => 
        counter_cry_Y(6), FCO => counter_cry_Z(6));
    
    \counter[15]\ : SLE
      port map(D => counter_s(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(15));
    
    \counter[29]\ : SLE
      port map(D => counter_s(29), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(29));
    
    \timestamp[8]\ : SLE
      port map(D => counter_Z(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(8));
    
    un1_prescaler_axbxc0 : CFG4
      generic map(INIT => x"33C4")

      port map(A => un6_enable_3_Z, B => counter_0_sqmuxa_0_Z, C
         => prescaler_Z(1), D => prescaler_Z(0), Y => 
        un1_prescaler_axbxc0_Z);
    
    un1_prescaler_ac0_1 : CFG4
      generic map(INIT => x"4000")

      port map(A => state_Z(0), B => enableTimestampGen, C => 
        prescaler_Z(1), D => prescaler_Z(0), Y => 
        un1_prescaler_c2);
    
    \prescaler[4]\ : SLE
      port map(D => prescaler_5_Z(4), CLK => sb_sb_0_FIC_0_CLK, 
        EN => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => prescaler_Z(4));
    
    \counter_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(11), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(10), S => counter_s(11), Y
         => counter_cry_Y(11), FCO => counter_cry_Z(11));
    
    \timestamp[2]\ : SLE
      port map(D => counter_Z(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(2));
    
    \counter_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(7), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(6), S => counter_s(7), Y => 
        counter_cry_Y(7), FCO => counter_cry_Z(7));
    
    \counter_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(1), C => \GND\, D => 
        \GND\, FCI => counter_s_830_FCO, S => counter_s(1), Y => 
        counter_cry_Y(1), FCO => counter_cry_Z(1));
    
    \counter[14]\ : SLE
      port map(D => counter_s(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(14));
    
    \timestamp[31]\ : SLE
      port map(D => counter_Z(31), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(31));
    
    state_0_sqmuxa : CFG2
      generic map(INIT => x"4")

      port map(A => state_Z(0), B => getTime, Y => 
        state_0_sqmuxa_Z);
    
    \timestamp[18]\ : SLE
      port map(D => counter_Z(18), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(18));
    
    \counter_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(12), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(11), S => counter_s(12), Y
         => counter_cry_Y(12), FCO => counter_cry_Z(12));
    
    \prescaler[1]\ : SLE
      port map(D => un1_prescaler_axbxc1_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        prescaler_Z(1));
    
    \counter_cry[30]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(30), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(29), S => counter_s(30), Y
         => counter_cry_Y(30), FCO => counter_cry_Z(30));
    
    \prescaler[2]\ : SLE
      port map(D => un1_prescaler_axbxc2_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        prescaler_Z(2));
    
    \counter[21]\ : SLE
      port map(D => counter_s(21), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(21));
    
    \timestamp[17]\ : SLE
      port map(D => counter_Z(17), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(17));
    
    \counter_cry[24]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(24), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(23), S => counter_s(24), Y
         => counter_cry_Y(24), FCO => counter_cry_Z(24));
    
    \counter[4]\ : SLE
      port map(D => counter_s(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(4));
    
    \timestamp[26]\ : SLE
      port map(D => counter_Z(26), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(26));
    
    \timestamp[15]\ : SLE
      port map(D => counter_Z(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(15));
    
    \counter[28]\ : SLE
      port map(D => counter_s(28), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(28));
    
    \timestamp[0]\ : SLE
      port map(D => counter_Z(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(0));
    
    \counter[5]\ : SLE
      port map(D => counter_s(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(5));
    
    \state[0]\ : SLE
      port map(D => state_0_sqmuxa_Z, CLK => sb_sb_0_FIC_0_CLK, 
        EN => enableTimestampGen, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        state_Z(0));
    
    \timestamp[5]\ : SLE
      port map(D => counter_Z(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(5));
    
    \counter_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(8), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(7), S => counter_s(8), Y => 
        counter_cry_Y(8), FCO => counter_cry_Z(8));
    
    \counter_cry[16]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(16), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(15), S => counter_s(16), Y
         => counter_cry_Y(16), FCO => counter_cry_Z(16));
    
    counter_s_830 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(0), C => \GND\, D => 
        \GND\, FCI => \VCC\, S => counter_s_830_S, Y => 
        counter_s_830_Y, FCO => counter_s_830_FCO);
    
    \counter_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(10), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(9), S => counter_s(10), Y => 
        counter_cry_Y(10), FCO => counter_cry_Z(10));
    
    \counter_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(5), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(4), S => counter_s(5), Y => 
        counter_cry_Y(5), FCO => counter_cry_Z(5));
    
    un1_prescaler_axbxc5 : CFG3
      generic map(INIT => x"78")

      port map(A => prescaler_Z(4), B => un1_prescaler_c4, C => 
        prescaler_Z(5), Y => un1_prescaler_axbxc5_Z);
    
    \counter_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(3), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(2), S => counter_s(3), Y => 
        counter_cry_Y(3), FCO => counter_cry_Z(3));
    
    \counter[31]\ : SLE
      port map(D => counter_s_Z(31), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(31));
    
    \timestamp[10]\ : SLE
      port map(D => counter_Z(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(10));
    
    \counter[12]\ : SLE
      port map(D => counter_s(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(12));
    
    \counter_cry[17]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(17), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(16), S => counter_s(17), Y
         => counter_cry_Y(17), FCO => counter_cry_Z(17));
    
    \counter_cry[29]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(29), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(28), S => counter_s(29), Y
         => counter_cry_Y(29), FCO => counter_cry_Z(29));
    
    \counter[1]\ : SLE
      port map(D => counter_s(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(1));
    
    \timestamp[23]\ : SLE
      port map(D => counter_Z(23), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(23));
    
    \timestamp[12]\ : SLE
      port map(D => counter_Z(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(12));
    
    \counter[3]\ : SLE
      port map(D => counter_s(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(3));
    
    \timestamp[21]\ : SLE
      port map(D => counter_Z(21), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(21));
    
    \counter[23]\ : SLE
      port map(D => counter_s(23), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(23));
    
    \counter[19]\ : SLE
      port map(D => counter_s(19), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(19));
    
    counter_0_sqmuxa_0 : CFG2
      generic map(INIT => x"4")

      port map(A => state_Z(0), B => enableTimestampGen, Y => 
        counter_0_sqmuxa_0_Z);
    
    \counter[20]\ : SLE
      port map(D => counter_s(20), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(20));
    
    un6_enable_3 : CFG4
      generic map(INIT => x"0040")

      port map(A => prescaler_Z(5), B => prescaler_Z(4), C => 
        prescaler_Z(3), D => prescaler_Z(2), Y => un6_enable_3_Z);
    
    \timestamp[29]\ : SLE
      port map(D => counter_Z(29), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(29));
    
    \counter_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(9), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(8), S => counter_s(9), Y => 
        counter_cry_Y(9), FCO => counter_cry_Z(9));
    
    counter_0_sqmuxa : CFG4
      generic map(INIT => x"0008")

      port map(A => un6_enable_3_Z, B => counter_0_sqmuxa_0_Z, C
         => prescaler_Z(1), D => prescaler_Z(0), Y => countere);
    
    \timestamp[3]\ : SLE
      port map(D => counter_Z(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(3));
    
    \timestamp[1]\ : SLE
      port map(D => counter_Z(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(1));
    
    GND_Z : GND
      port map(Y => \GND\);
    
    \counter_cry[28]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(28), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(27), S => counter_s(28), Y
         => counter_cry_Y(28), FCO => counter_cry_Z(28));
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    \counter[27]\ : SLE
      port map(D => counter_s(27), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(27));
    
    \counter[11]\ : SLE
      port map(D => counter_s(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(11));
    
    \timestamp[30]\ : SLE
      port map(D => counter_Z(30), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(30));
    
    prescaler_2_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => state_Z(0), B => enableTimestampGen, Y => 
        prescaler_2_sqmuxa_Z);
    
    \counter[30]\ : SLE
      port map(D => counter_s(30), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(30));
    
    \counter[18]\ : SLE
      port map(D => counter_s(18), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(18));
    
    \prescaler[3]\ : SLE
      port map(D => prescaler_5_Z(3), CLK => sb_sb_0_FIC_0_CLK, 
        EN => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => prescaler_Z(3));
    
    \counter_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(2), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(1), S => counter_s(2), Y => 
        counter_cry_Y(2), FCO => counter_cry_Z(2));
    
    \counter_cry[14]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(14), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(13), S => counter_s(14), Y
         => counter_cry_Y(14), FCO => counter_cry_Z(14));
    
    \timestamp[14]\ : SLE
      port map(D => counter_Z(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(14));
    
    \counter_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(4), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(3), S => counter_s(4), Y => 
        counter_cry_Y(4), FCO => counter_cry_Z(4));
    
    \counter_cry[25]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(25), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(24), S => counter_s(25), Y
         => counter_cry_Y(25), FCO => counter_cry_Z(25));
    
    \timestamp[28]\ : SLE
      port map(D => counter_Z(28), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(28));
    
    \counter_cry[23]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(23), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(22), S => counter_s(23), Y
         => counter_cry_Y(23), FCO => counter_cry_Z(23));
    
    \prescaler_5[4]\ : CFG3
      generic map(INIT => x"12")

      port map(A => un1_prescaler_c4, B => countere, C => 
        prescaler_Z(4), Y => prescaler_5_Z(4));
    
    \timestamp[27]\ : SLE
      port map(D => counter_Z(27), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(27));
    
    \timestamp[25]\ : SLE
      port map(D => counter_Z(25), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(25));
    
    \timestamp[9]\ : SLE
      port map(D => counter_Z(9), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(9));
    
    \counter_cry[19]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => counter_Z(19), C => \GND\, D => 
        \GND\, FCI => counter_cry_Z(18), S => counter_s(19), Y
         => counter_cry_Y(19), FCO => counter_cry_Z(19));
    
    \counter[26]\ : SLE
      port map(D => counter_s(26), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(26));
    
    \counter[13]\ : SLE
      port map(D => counter_s(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(13));
    
    \counter[0]\ : SLE
      port map(D => counter_s(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(0));
    
    \timestamp[6]\ : SLE
      port map(D => counter_Z(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => prescaler_2_sqmuxa_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        TimeStampValue(6));
    
    \counter[10]\ : SLE
      port map(D => counter_s(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(10));
    
    \counter[9]\ : SLE
      port map(D => counter_s(9), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(9));
    
    \counter[25]\ : SLE
      port map(D => counter_s(25), CLK => sb_sb_0_FIC_0_CLK, EN
         => countere, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(25));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Memory is

    port( sb_sb_0_STAMP_PADDR   : in    std_logic_vector(11 downto 0);
          dataReady_0           : in    std_logic;
          STAMP_0_data_frame    : in    std_logic_vector(63 downto 0);
          sb_sb_0_Memory_PRDATA : out   std_logic_vector(31 downto 0);
          sb_sb_0_STAMP_PWDATA  : in    std_logic_vector(31 downto 0);
          nCS1_c                : out   std_logic;
          nCS2_c                : out   std_logic;
          MISO_c                : in    std_logic;
          SCLK_c                : out   std_logic;
          mosi_1                : out   std_logic;
          mosi_cl               : out   std_logic;
          sb_sb_0_STAMP_PENABLE : in    std_logic;
          sb_sb_0_STAMP_PWRITE  : in    std_logic;
          sb_sb_0_Memory_PSELx  : in    std_logic;
          un1_APBState_1_5_1z   : out   std_logic;
          resetn                : in    std_logic;
          sb_sb_0_Memory_PREADY : out   std_logic;
          GPIO_6_M2F_c          : in    std_logic;
          sb_sb_0_FIC_0_CLK     : in    std_logic;
          resetn_arst           : in    std_logic
        );

end Memory;

architecture DEF_ARCH of Memory is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component spi_master_2_32
    port( SPITransmitReg    : in    std_logic_vector(31 downto 0) := (others => 'U');
          SPIaddr_0         : in    std_logic := 'U';
          SPIRecReg         : out   std_logic_vector(31 downto 0);
          enable            : in    std_logic := 'U';
          InternalBusy      : out   std_logic;
          mosi_cl_1z        : out   std_logic;
          mosi_1_1z         : out   std_logic;
          resetn            : in    std_logic := 'U';
          SCLK_c            : out   std_logic;
          MISO_c            : in    std_logic := 'U';
          nCS2_c            : out   std_logic;
          resetn_arst       : in    std_logic := 'U';
          nCS1_c            : out   std_logic;
          sb_sb_0_FIC_0_CLK : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component ram
    port( InternalData2Memory : in    std_logic_vector(31 downto 0) := (others => 'U');
          InternalAddr2Memory : in    std_logic_vector(8 downto 0) := (others => 'U');
          InternalDataFromMem : out   std_logic_vector(31 downto 0);
          resetn              : in    std_logic := 'U';
          WriteEnable         : in    std_logic := 'U';
          sb_sb_0_FIC_0_CLK   : in    std_logic := 'U';
          resetn_arst         : in    std_logic := 'U'
        );
  end component;

  component Timestamp
    port( TimeStampValue     : out   std_logic_vector(31 downto 0);
          getTime            : in    std_logic := 'U';
          enableTimestampGen : in    std_logic := 'U';
          sb_sb_0_FIC_0_CLK  : in    std_logic := 'U';
          resetn_arst        : in    std_logic := 'U'
        );
  end component;

    signal \un1_APBState_1_5_1z\ : std_logic;
    signal ControllUnitState_RNI2VHT_Z : 
        std_logic_vector(14 to 14);
    signal counter_Z : std_logic_vector(1 downto 0);
    signal ConfigStatusReg_Z : std_logic_vector(31 downto 0);
    signal MemoryPageSize : std_logic_vector(15 downto 0);
    signal ConfigStatusReg_40 : std_logic_vector(29 to 29);
    signal ConfigStatusReg_26 : std_logic_vector(30 to 30);
    signal StartAddrReg_Z : std_logic_vector(31 downto 0);
    signal readmemorycounter_Z : std_logic_vector(3 downto 0);
    signal readmemorycounter_6 : std_logic_vector(1 to 1);
    signal pageaddr : std_logic_vector(30 downto 0);
    signal pageaddr_5_i_m4 : std_logic_vector(30 downto 0);
    signal pageaddr_5 : std_logic_vector(27 to 27);
    signal CurrentAddrReg_Z : std_logic_vector(31 downto 0);
    signal StampFSMPC_Z : std_logic_vector(8 downto 0);
    signal StampFSMPC_6 : std_logic_vector(8 downto 2);
    signal PRDATA_8 : std_logic_vector(31 downto 0);
    signal StampFSMPC_6_Z : std_logic_vector(1 to 1);
    signal InternalData2Memory_Z : std_logic_vector(31 downto 0);
    signal InternalData2Memory_27 : 
        std_logic_vector(31 downto 0);
    signal Command_Z : std_logic_vector(7 downto 0);
    signal SPITransmitReg_Z : std_logic_vector(31 downto 0);
    signal SPITransmitReg_13 : std_logic_vector(31 downto 0);
    signal tempcounter_Z : std_logic_vector(8 downto 0);
    signal tempcounter_7_iv_i : std_logic_vector(7 downto 0);
    signal tempcounter_7 : std_logic_vector(1 to 1);
    signal InternalAddr2Memory_Z : std_logic_vector(8 downto 0);
    signal InternalAddr2Memory_34 : std_logic_vector(8 downto 0);
    signal Stamp1ShadowReg1_Z : std_logic_vector(31 downto 0);
    signal Stamp1ShadowReg2_Z : std_logic_vector(31 downto 0);
    signal ReadMemoryShadowReg_Z : std_logic_vector(31 downto 0);
    signal InternalDataFromMem : std_logic_vector(31 downto 0);
    signal CommandReg_Z : std_logic_vector(31 downto 0);
    signal readmemorylimitedcnt_Z : std_logic_vector(8 downto 0);
    signal readmemorylimitedcnt_5 : std_logic_vector(8 downto 0);
    signal readmemoryaddrcounter_Z : 
        std_logic_vector(31 downto 23);
    signal readmemoryaddrcounter_3_Z : 
        std_logic_vector(8 downto 0);
    signal memorycnt_Z : std_logic_vector(8 downto 1);
    signal memorycnt_6 : std_logic_vector(8 downto 2);
    signal MemoryPageSize_Z : std_logic_vector(13 downto 2);
    signal ControllUnitState_Z : std_logic_vector(14 downto 0);
    signal ControllUnitState_ns : std_logic_vector(13 downto 0);
    signal ControllUnitSubState_Z : std_logic_vector(1 downto 0);
    signal ControllUnitSubState_ns : std_logic_vector(0 to 0);
    signal SPIaddr_Z : std_logic_vector(0 to 0);
    signal SPIaddr_15 : std_logic_vector(0 to 0);
    signal isfirstrun_Z : std_logic_vector(0 to 0);
    signal ReadMemoryState_Z : std_logic_vector(8 downto 0);
    signal ReadMemoryState_ns_i_i_Z : std_logic_vector(8 to 8);
    signal APBState_Z : std_logic_vector(1 downto 0);
    signal APBState_ns : std_logic_vector(1 downto 0);
    signal ReadMemoryState_ns : std_logic_vector(5 downto 4);
    signal APB3ReadMemoryLimitedState_Z : 
        std_logic_vector(5 downto 0);
    signal APB3ReadMemoryLimitedState_ns : 
        std_logic_vector(4 downto 0);
    signal APB3ReadMemoryLimitedState_RNI12J4_Y : 
        std_logic_vector(5 to 5);
    signal SPIState_Z : std_logic_vector(4 downto 0);
    signal SPIState_ns : std_logic_vector(3 to 3);
    signal APB3ReadMemoryLimitedState_RNI12J4_S : 
        std_logic_vector(5 to 5);
    signal readmemorylimitedcnt_RNI1LOJ_S : 
        std_logic_vector(0 to 0);
    signal readmemorylimitedcnt_RNI1LOJ_Y : 
        std_logic_vector(0 to 0);
    signal readmemorylimitedcnt_RNI29U21_S : 
        std_logic_vector(1 to 1);
    signal readmemorylimitedcnt_RNI29U21_Y : 
        std_logic_vector(1 to 1);
    signal readmemorylimitedcnt_RNI4U3I1_S : 
        std_logic_vector(2 to 2);
    signal readmemorylimitedcnt_RNI4U3I1_Y : 
        std_logic_vector(2 to 2);
    signal readmemorylimitedcnt_RNI7K912_S : 
        std_logic_vector(3 to 3);
    signal readmemorylimitedcnt_RNI7K912_Y : 
        std_logic_vector(3 to 3);
    signal readmemorylimitedcnt_RNIBBFG2_S : 
        std_logic_vector(4 to 4);
    signal readmemorylimitedcnt_RNIBBFG2_Y : 
        std_logic_vector(4 to 4);
    signal readmemorylimitedcnt_RNIG3LV2_S : 
        std_logic_vector(5 to 5);
    signal readmemorylimitedcnt_RNIG3LV2_Y : 
        std_logic_vector(5 to 5);
    signal readmemorylimitedcnt_RNIMSQE3_S : 
        std_logic_vector(6 to 6);
    signal readmemorylimitedcnt_RNIMSQE3_Y : 
        std_logic_vector(6 to 6);
    signal readmemorylimitedcnt_5_RNO_FCO : 
        std_logic_vector(8 to 8);
    signal readmemorylimitedcnt_5_RNO_S : 
        std_logic_vector(8 to 8);
    signal readmemorylimitedcnt_5_RNO_Y : 
        std_logic_vector(8 to 8);
    signal readmemorylimitedcnt_RNITM0U3_S : 
        std_logic_vector(7 to 7);
    signal readmemorylimitedcnt_RNITM0U3_Y : 
        std_logic_vector(7 to 7);
    signal un23_0_0_Z : std_logic_vector(2 to 2);
    signal un23_0_a2_1_0_Z : std_logic_vector(2 to 2);
    signal un23_1_Z : std_logic_vector(1 to 1);
    signal un23_a3_0 : std_logic_vector(1 to 1);
    signal TimeStampValue : std_logic_vector(31 downto 0);
    signal InternalAddr2Memory_34_m2_1_1 : 
        std_logic_vector(1 downto 0);
    signal SPIState_RNO_1_Z : std_logic_vector(2 to 2);
    signal SPITransmitReg_RNO_1_Z : std_logic_vector(4 downto 0);
    signal SPIState_RNO_5_Z : std_logic_vector(2 to 2);
    signal ConfigStatusReg_26_0_m2_1 : 
        std_logic_vector(30 to 30);
    signal ConfigStatusReg_26_0_1 : std_logic_vector(30 to 30);
    signal ConfigStatusReg_26_0_a2_1 : 
        std_logic_vector(30 to 30);
    signal InternalAddr2Memory_34_m2 : 
        std_logic_vector(8 downto 0);
    signal InternalAddr2Memory_34_m2_1_0 : 
        std_logic_vector(8 to 8);
    signal InternalAddr2Memory_34_1 : 
        std_logic_vector(7 downto 2);
    signal InternalAddr2Memory_34_m0 : 
        std_logic_vector(7 downto 2);
    signal InternalAddr2Memory_34_m4 : std_logic_vector(1 to 1);
    signal SPIRecReg : std_logic_vector(31 downto 0);
    signal InternalData2Memory_27_0_iv_0_0 : 
        std_logic_vector(31 downto 0);
    signal InternalData2Memory_27_0_iv_0 : 
        std_logic_vector(30 downto 11);
    signal ControllUnitSubState_ns_i_a7_0_3_Z : 
        std_logic_vector(1 to 1);
    signal ControllUnitSubState_ns_i_a7_0_2_Z : 
        std_logic_vector(1 to 1);
    signal ControllUnitSubState_ns_0_0_a2_1_Z : 
        std_logic_vector(0 to 0);
    signal ControllUnitState_ns_i_0_a2_1 : 
        std_logic_vector(14 to 14);
    signal ControllUnitSubState_ns_i_a7_4_4_Z : 
        std_logic_vector(1 to 1);
    signal ControllUnitSubState_ns_i_a7_4_3_Z : 
        std_logic_vector(1 to 1);
    signal ControllUnitState_ns_i_a2_3_Z : 
        std_logic_vector(11 to 11);
    signal ReadMemoryState_ns_i_0_a3_2_7_Z : 
        std_logic_vector(3 to 3);
    signal ReadMemoryState_ns_i_0_a3_2_6_Z : 
        std_logic_vector(3 to 3);
    signal ControllUnitSubState_ns_i_a7_0_Z : 
        std_logic_vector(1 to 1);
    signal ReadMemoryState_ns_i_o4_3_Z : 
        std_logic_vector(0 to 0);
    signal ConfigStatusReg_RNO_2_Z : std_logic_vector(4 to 4);
    signal pageaddr_m : std_logic_vector(1 to 1);
    signal SPIState_RNI27U44_Z : std_logic_vector(1 to 1);
    signal InternalData2Memory_27_0_iv_0_1 : 
        std_logic_vector(28 downto 0);
    signal InternalData2Memory_27_0_iv_1 : 
        std_logic_vector(25 downto 11);
    signal ControllUnitSubState_ns_i_0_Z : 
        std_logic_vector(1 to 1);
    signal ControllUnitSubState_ns_i_a7_4_5_Z : 
        std_logic_vector(1 to 1);
    signal ReadMemoryState_ns_i_0_a3_2_8_Z : 
        std_logic_vector(3 to 3);
    signal ControllUnitState_ns_i_0_1_Z : 
        std_logic_vector(11 to 11);
    signal InternalAddr2Memory_34_m5 : 
        std_logic_vector(8 downto 0);
    signal PRDATA_8_0_iv_0_3 : std_logic_vector(31 downto 0);
    signal PRDATA_8_0_iv_0_2 : std_logic_vector(31 downto 0);
    signal PRDATA_8_0_iv_0_1 : std_logic_vector(31 downto 0);
    signal PRDATA_8_0_iv_0_0 : std_logic_vector(31 downto 0);
    signal InternalData2Memory_27_0_iv_0_3 : 
        std_logic_vector(28 downto 0);
    signal InternalData2Memory_27_0_iv_3 : 
        std_logic_vector(25 downto 11);
    signal InternalData2Memory_27_0_iv_2 : 
        std_logic_vector(30 downto 24);
    signal InternalData2Memory_27_0_iv_0_2 : 
        std_logic_vector(31 to 31);
    signal ControllUnitSubState_ns_i_1_Z : 
        std_logic_vector(1 to 1);
    signal ControllUnitState_ns_i_0_a2_0_1_Z : 
        std_logic_vector(14 to 14);
    signal ControllUnitState_ns_i_0_2_Z : 
        std_logic_vector(11 to 11);
    signal ControllUnitSubState_ns_i_2_Z : 
        std_logic_vector(1 to 1);
    signal ReadMemoryState_ns_i_0_0_Z : std_logic_vector(3 to 3);
    signal PRDATA_8_0_iv_0_6 : std_logic_vector(31 downto 0);
    signal ControllUnitState_ns_i_0_0_Z : 
        std_logic_vector(14 to 14);
    signal N_1541_i, \VCC\, N_140_mux_i, \GND\, N_4253_i, 
        N_4340_i, N_249_i, N_88, N_87, N_85_i, N_252_i, 
        StartAddrReg_0_sqmuxa, N_4260_i, N_4261_i, N_4262_i, 
        N_4371, N_4370, N_4369, un1_currentaddrreg_cry_28_S, 
        N_4294_i, un1_currentaddrreg_cry_29_S, 
        un1_currentaddrreg_cry_30_S, un1_currentaddrreg_cry_30_Z, 
        un1_currentaddrreg_cry_13_S, un1_currentaddrreg_cry_14_S, 
        un1_currentaddrreg_cry_15_S, un1_currentaddrreg_cry_16_S, 
        un1_currentaddrreg_cry_17_S, un1_currentaddrreg_cry_18_S, 
        un1_currentaddrreg_cry_19_S, un1_currentaddrreg_cry_20_S, 
        un1_currentaddrreg_cry_21_S, un1_currentaddrreg_cry_22_S, 
        un1_currentaddrreg_cry_23_S, un1_currentaddrreg_cry_24_S, 
        un1_currentaddrreg_cry_25_S, un1_currentaddrreg_cry_26_S, 
        un1_currentaddrreg_cry_27_S, N_1246_i, 
        un1_currentaddrreg_cry_0_Y, un1_currentaddrreg_cry_1_S, 
        un1_currentaddrreg_cry_2_S, un1_currentaddrreg_cry_3_S, 
        un1_currentaddrreg_cry_4_S, un1_currentaddrreg_cry_5_S, 
        un1_currentaddrreg_cry_6_S, un1_currentaddrreg_cry_7_S, 
        un1_currentaddrreg_cry_8_S, un1_currentaddrreg_cry_9_S, 
        un1_currentaddrreg_cry_10_S, un1_currentaddrreg_cry_11_S, 
        un1_currentaddrreg_cry_12_S, un1_APBState_1_i, N_746_i, 
        InternalData2Memory_0_sqmuxa_6_i_Z, N_172_i, 
        Command_1_sqmuxa_1_i_Z, N_170_i, N_168_i, N_166_i, N_16, 
        un1_enabletimestampgen2_1_i, N_139_i, N_4295_i, N_4296_i, 
        N_4297_i, N_4298_i, N_4299_i, N_180_i, N_178_i, N_176_i, 
        N_174_i, InternalAddr2Memory_0_sqmuxa_i_Z, N_1080_i, 
        ReadMemoryShadowReg_0_sqmuxa_i_Z, Command_1_sqmuxa, 
        un1_readmemoryaddrcounter_cry_1_S, 
        un1_readmemoryaddrcounter_cry_2_S, 
        un1_readmemoryaddrcounter_cry_3_S, 
        un1_readmemoryaddrcounter_cry_4_S, 
        un1_readmemoryaddrcounter_cry_5_S, 
        un1_readmemoryaddrcounter_cry_6_S, memorycnt_6_cry_0_0_Y, 
        N_2624_2, N_161, N_7_0, N_2629_i, N_127, enable, 
        un1_SPIState_8, enableSPI_0_sqmuxa_3_i_Z, getTime_Z, 
        getTime_3, WriteEnable_Z, N_4265_i, 
        WriteEnable_0_sqmuxa_i_Z, isfirstrun_1_sqmuxa, N_1539_i, 
        N_2554_i, N_2550_i, N_2471_i, N_44, N_2475_i, N_2477_i, 
        N_101, N_145_mux, N_154_mux_i, N_157_mux, N_70, N_42_0, 
        enableTimestampGen_Z, un1_readmemorylimitedcnt_cry_0_cy, 
        un1_readmemorylimitedcnt_cry_0, 
        un1_readmemorylimitedcnt_cry_1, 
        un1_readmemorylimitedcnt_cry_2, 
        un1_readmemorylimitedcnt_cry_3, 
        un1_readmemorylimitedcnt_cry_4, 
        un1_readmemorylimitedcnt_cry_5, 
        un1_readmemorylimitedcnt_cry_6, 
        un1_readmemorylimitedcnt_cry_7, memorycnt_6_cry_0, 
        memorycnt_6_cry_0_0_S, N_1255_i, memorycnt_6_cry_1, 
        memorycnt_6_cry_1_0_Y, memorycnt_6_cry_2, 
        memorycnt_6_cry_2_0_Y, memorycnt_6_cry_3, 
        memorycnt_6_cry_3_Y, memorycnt_6_cry_4, 
        memorycnt_6_cry_4_Y, memorycnt_6_cry_5, 
        memorycnt_6_cry_5_Y, memorycnt_6_s_7_FCO, 
        memorycnt_6_s_7_Y, memorycnt_6_cry_6, memorycnt_6_cry_6_Y, 
        un1_memorycnt_1_cry_1_Z, un1_memorycnt_1_cry_1_S, 
        un1_memorycnt_1_cry_1_Y, N_1260, un1_memorycnt_1_cry_2_Z, 
        un1_memorycnt_1_cry_2_S, un1_memorycnt_1_cry_2_Y, N_1262, 
        un1_memorycnt_1_cry_3_Z, un1_memorycnt_1_cry_3_S, 
        un1_memorycnt_1_cry_3_Y, N_761, N_762, N_4343, 
        un1_memorycnt_1_cry_4_Z, un1_memorycnt_1_cry_4_S, 
        un1_memorycnt_1_cry_4_Y, un1_memorycnt_1_cry_5_Z, 
        un1_memorycnt_1_cry_5_S, un1_memorycnt_1_cry_5_Y, 
        un1_memorycnt_1_cry_6_Z, un1_memorycnt_1_cry_6_S, 
        un1_memorycnt_1_cry_6_Y, un1_memorycnt_1_s_8_FCO, 
        un1_memorycnt_1_s_8_S, un1_memorycnt_1_s_8_Y, 
        un1_memorycnt_1_cry_7_Z, un1_memorycnt_1_cry_7_S, 
        un1_memorycnt_1_cry_7_Y, un1_currentaddrreg_cry_0_Z, 
        un1_currentaddrreg_cry_0_S, un1_currentaddrreg_cry_1_Z, 
        un1_currentaddrreg_cry_1_Y, un1_currentaddrreg_cry_2_Z, 
        un1_currentaddrreg_cry_2_Y, un1_currentaddrreg_cry_3_Z, 
        un1_currentaddrreg_cry_3_Y, un1_currentaddrreg_cry_4_Z, 
        un1_currentaddrreg_cry_4_Y, un1_currentaddrreg_cry_5_Z, 
        un1_currentaddrreg_cry_5_Y, un1_currentaddrreg_cry_6_Z, 
        un1_currentaddrreg_cry_6_Y, un1_currentaddrreg_cry_7_Z, 
        un1_currentaddrreg_cry_7_Y, un1_currentaddrreg_cry_8_Z, 
        un1_currentaddrreg_cry_8_Y, un1_currentaddrreg_cry_9_Z, 
        un1_currentaddrreg_cry_9_Y, un1_currentaddrreg_cry_10_Z, 
        un1_currentaddrreg_cry_10_Y, un1_currentaddrreg_cry_11_Z, 
        un1_currentaddrreg_cry_11_Y, un1_currentaddrreg_cry_12_Z, 
        un1_currentaddrreg_cry_12_Y, un1_currentaddrreg_cry_13_Z, 
        un1_currentaddrreg_cry_13_Y, un1_currentaddrreg_cry_14_Z, 
        un1_currentaddrreg_cry_14_Y, un1_currentaddrreg_cry_15_Z, 
        un1_currentaddrreg_cry_15_Y, un1_currentaddrreg_cry_16_Z, 
        un1_currentaddrreg_cry_16_Y, un1_currentaddrreg_cry_17_Z, 
        un1_currentaddrreg_cry_17_Y, un1_currentaddrreg_cry_18_Z, 
        un1_currentaddrreg_cry_18_Y, un1_currentaddrreg_cry_19_Z, 
        un1_currentaddrreg_cry_19_Y, un1_currentaddrreg_cry_20_Z, 
        un1_currentaddrreg_cry_20_Y, un1_currentaddrreg_cry_21_Z, 
        un1_currentaddrreg_cry_21_Y, un1_currentaddrreg_cry_22_Z, 
        un1_currentaddrreg_cry_22_Y, un1_currentaddrreg_cry_23_Z, 
        un1_currentaddrreg_cry_23_Y, un1_currentaddrreg_cry_24_Z, 
        un1_currentaddrreg_cry_24_Y, un1_currentaddrreg_cry_25_Z, 
        un1_currentaddrreg_cry_25_Y, un1_currentaddrreg_cry_26_Z, 
        un1_currentaddrreg_cry_26_Y, un1_currentaddrreg_cry_27_Z, 
        un1_currentaddrreg_cry_27_Y, un1_currentaddrreg_cry_28_Z, 
        un1_currentaddrreg_cry_28_Y, un1_currentaddrreg_cry_29_Z, 
        un1_currentaddrreg_cry_29_Y, un1_currentaddrreg_cry_30_Y, 
        un8_tempcounter_s_1_835_FCO, un8_tempcounter_s_1_835_S, 
        un8_tempcounter_s_1_835_Y, un8_tempcounter_cry_1_Z, 
        un8_tempcounter_cry_1_S, un8_tempcounter_cry_1_Y, 
        un8_tempcounter_cry_2_Z, un8_tempcounter_cry_2_S, 
        un8_tempcounter_cry_2_Y, un8_tempcounter_cry_3_Z, 
        un8_tempcounter_cry_3_S, un8_tempcounter_cry_3_Y, 
        un8_tempcounter_cry_4_Z, un8_tempcounter_cry_4_S, 
        un8_tempcounter_cry_4_Y, un8_tempcounter_cry_5_Z, 
        un8_tempcounter_cry_5_S, un8_tempcounter_cry_5_Y, 
        un8_tempcounter_cry_6_Z, un8_tempcounter_cry_6_S, 
        un8_tempcounter_cry_6_Y, un8_tempcounter_s_8_FCO, 
        un8_tempcounter_s_8_S, un8_tempcounter_s_8_Y, 
        un8_tempcounter_cry_7_Z, un8_tempcounter_cry_7_S, 
        un8_tempcounter_cry_7_Y, 
        un1_readmemoryaddrcounter_s_0_836_FCO, 
        un1_readmemoryaddrcounter_s_0_836_S, 
        un1_readmemoryaddrcounter_s_0_836_Y, 
        un1_readmemoryaddrcounter_cry_0_Z, 
        un1_readmemoryaddrcounter_cry_0_S, 
        un1_readmemoryaddrcounter_cry_0_Y, 
        un1_readmemoryaddrcounter_cry_1_Z, 
        un1_readmemoryaddrcounter_cry_1_Y, 
        un1_readmemoryaddrcounter_cry_2_Z, 
        un1_readmemoryaddrcounter_cry_2_Y, 
        un1_readmemoryaddrcounter_cry_3_Z, 
        un1_readmemoryaddrcounter_cry_3_Y, 
        un1_readmemoryaddrcounter_cry_4_Z, 
        un1_readmemoryaddrcounter_cry_4_Y, 
        un1_readmemoryaddrcounter_cry_5_Z, 
        un1_readmemoryaddrcounter_cry_5_Y, 
        un1_readmemoryaddrcounter_cry_6_Z, 
        un1_readmemoryaddrcounter_cry_6_Y, 
        un1_readmemoryaddrcounter_s_8_FCO, 
        un1_readmemoryaddrcounter_s_8_S, 
        un1_readmemoryaddrcounter_s_8_Y, 
        un1_readmemoryaddrcounter_cry_7_Z, 
        un1_readmemoryaddrcounter_cry_7_S, 
        un1_readmemoryaddrcounter_cry_7_Y, SPIaddr_0_sqmuxa_3, 
        N_23_0, SPIaddr_3_sqmuxa_1, N_4343_i, N_1232_i, N_4527, 
        N_138, N_143_mux, m41_0_1, m41_0_2_1, SPIState_1_sqmuxa, 
        SPIState_m2_e_1_0_Z, SPIState_m2_e_1, SPIState_m2_e_1_1_Z, 
        N_4272_i, N_4270, N_13_mux_1, N_54, N_13_mux_0, N_13_mux, 
        N_1034, N_4_23, N_15_mux_22, N_4_22, N_15_mux_21, N_4_21, 
        N_15_mux_20, N_4_20, N_15_mux_19, N_4_19, N_15_mux_18, 
        N_4_18, N_15_mux_17, N_4_17, N_15_mux_16, N_4_16, 
        N_15_mux_15, N_4_15, N_15_mux_14, N_4_14, N_15_mux_13, 
        N_4_13, N_15_mux_12, N_4_12, N_15_mux_11, N_4_11, 
        N_15_mux_10, N_4_10, N_15_mux_9, N_4_9, N_15_mux_8, N_4_8, 
        N_15_mux_7, N_4_7, N_15_mux_6, N_4_6, N_15_mux_5, N_4_5, 
        N_15_mux_4, N_4_4, N_15_mux_3, N_4_3, N_15_mux_2, N_4_2, 
        N_15_mux_1, N_4_1, N_15_mux_0, N_4_0, N_15_mux, m33_e_0, 
        counter9, m46_1_1_0, m46_0, m46_1_1, N_4340, N_2624, 
        m98_xx_mm_1, N_149_mux, N_2471_i_1, N_2496, N_4274, N_68, 
        N_62, N_154_mux_i_1_0, N_21_0, m46_1_1_0_1, m46_1_1_tz, 
        N_1316_i, N_4354, InternalAddr2Memory_34_sm0, m94_1_1, 
        N_89, N_146, N_2496_i, m87_0_1, m87_m7_0, r_N_6_mux, 
        m84_m7_0, m86_0_1, m86_m7_0, N_19_0, m106_1_1, 
        InternalAddr2Memory_34_2, InternalAddr2Memory_34_6, 
        InternalAddr2Memory_34_10, InternalAddr2Memory_34_14, 
        InternalAddr2Memory_34_18, InternalAddr2Memory_34_22, 
        m84_N_13_mux, d_N_5_mux, N_765_1, N_1261_i, 
        ConfigStatusReg_24_sn_N_5, N_81, N_4268, N_1254, N_4344, 
        InternalData2Memory_3_sqmuxa_Z, N_1128, N_4351, 
        enableSPI_1_sqmuxa_1_0_Z, N_1257_i, N_2648, N_4342, 
        N_1041, N_4339, N_2624_1, N_4258, N_4423, N_155_mux_i, 
        N_4358, PRDATA_17_sqmuxa_2_Z, m73_m2_e_0_0, 
        Command_1_sqmuxa_0_a2_1_0_Z, un1_APBState_1_1_Z, 
        un1_enabletimestampgen2_5_6_Z, 
        un1_enabletimestampgen2_5_3_Z, 
        un1_enabletimestampgen2_5_2_Z, 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_1_Z, m60_e_5, m60_e_4, 
        ControllUnitState_tr25_0_a2_5_Z, 
        ControllUnitState_tr25_0_a2_4_Z, m17_e_1, N_1298, N_2631, 
        un1_paddr_3, N_1302, N_1035, InternalBusy, 
        un1_SPIState_8_0_a3_0_Z, InternalData2Memory_5_sqmuxa_Z, 
        N_712, N_144, InternalData2Memory_4_sqmuxa_Z, 
        un1_APBState_1_2_0_Z, N_4535, un1_ControllUnitState_9, 
        PRDATA_17_sqmuxa_8_Z, N_1025, N_1026, N_1028, N_1029, 
        N_1031, N_1032, N_4335, N_1045, N_1030, N_4546, N_4266, 
        N_4424, N_4348, N_4347, MemoryPageSize_1_sqmuxa_0_o4_0_Z, 
        m73_m2_e_1, m84_m7_1, un1_enabletimestampgen2_5_8_Z, 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_7_Z, 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_6_Z, 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_2_Z, 
        un1_enabletimestampgen2_7_0_0_Z, N_1185, 
        Command_1_sqmuxa_0_a2_0_Z, N_4350, N_1508_i, N_1033, 
        N_4547, ConfigStatusReg_24_sn_N_11_mux, m73_m2_e_2, 
        un1_enabletimestampgen2_5_7_Z, N_1186, N_5700, 
        PRDATA_17_sqmuxa_Z, N_139_mux, N_4614, N_4346, 
        un1_enableSPI_1_sqmuxa_1_i, N_4259, N_95, N_4349, 
        N_4254_i, enableSPI_0_sqmuxa_2, 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_8_Z, N_765, N_80, 
        N_4286, N_734, N_4353, N_102, N_50_0, N_2641, N_71, 
        N_31_0, N_150_mux, N_327, N_1514, N_1513, N_1512, N_1329, 
        N_1328, N_1327, N_1326, N_1325, N_1324, N_1323, N_1322, 
        N_1321, N_886, N_885, N_884, N_883, N_882, N_881, N_880, 
        N_879, N_878, N_877, N_876, N_875, N_874, N_873, N_872, 
        N_794, N_793, N_792, N_732, N_731, N_730, N_729, N_728, 
        N_727, N_655, N_654, N_653, N_652, N_651, N_322
         : std_logic;

    for all : spi_master_2_32
	Use entity work.spi_master_2_32(DEF_ARCH);
    for all : ram
	Use entity work.ram(DEF_ARCH);
    for all : Timestamp
	Use entity work.Timestamp(DEF_ARCH);
begin 

    un1_APBState_1_5_1z <= \un1_APBState_1_5_1z\;

    enableSPI_0_sqmuxa_3_i : CFG4
      generic map(INIT => x"DDD5")

      port map(A => enableSPI_0_sqmuxa_2, B => GPIO_6_M2F_c, C
         => ControllUnitState_Z(1), D => enableSPI_1_sqmuxa_1_0_Z, 
        Y => enableSPI_0_sqmuxa_3_i_Z);
    
    \Command_RNO[7]\ : CFG2
      generic map(INIT => x"4")

      port map(A => SPIState_RNI27U44_Z(1), B => 
        sb_sb_0_STAMP_PWDATA(31), Y => N_166_i);
    
    \mainProcess.pageaddr_5_i_m4[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(3), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(3), Y => pageaddr_5_i_m4(3));
    
    \SPITransmitReg[8]\ : SLE
      port map(D => SPITransmitReg_13(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(8));
    
    \StampFSMR1[4]\ : SLE
      port map(D => pageaddr_5_i_m4(4), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(4));
    
    \SPITransmitReg_RNO[25]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_6, B => InternalDataFromMem(25), C => 
        N_54, D => N_15_mux_5, Y => SPITransmitReg_13(25));
    
    \readmemorylimitedcnt_RNIG3LV2[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemorylimitedcnt_Z(5), C => 
        \GND\, D => \GND\, FCI => un1_readmemorylimitedcnt_cry_4, 
        S => readmemorylimitedcnt_RNIG3LV2_S(5), Y => 
        readmemorylimitedcnt_RNIG3LV2_Y(5), FCO => 
        un1_readmemorylimitedcnt_cry_5);
    
    \CommandReg[4]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(4));
    
    \mainProcess.PRDATA_8_0_iv_0_a2_10[12]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => sb_sb_0_STAMP_PADDR(2), B => 
        sb_sb_0_STAMP_PADDR(5), C => sb_sb_0_STAMP_PADDR(4), D
         => sb_sb_0_STAMP_PADDR(3), Y => N_1032);
    
    un1_currentaddrreg_cry_30 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(30), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_29_Z, S => 
        un1_currentaddrreg_cry_30_S, Y => 
        un1_currentaddrreg_cry_30_Y, FCO => 
        un1_currentaddrreg_cry_30_Z);
    
    SPIState_1_sqmuxa_0_a2_0 : CFG4
      generic map(INIT => x"8000")

      port map(A => sb_sb_0_STAMP_PADDR(2), B => 
        sb_sb_0_STAMP_PADDR(5), C => sb_sb_0_STAMP_PADDR(4), D
         => sb_sb_0_STAMP_PADDR(3), Y => N_1026);
    
    \SPIaddr[0]\ : SLE
      port map(D => SPIaddr_15(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_127, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => SPIaddr_Z(0));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[17]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(17), B => 
        TimeStampValue(17), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(17));
    
    \readmemoryaddrcounter[29]\ : SLE
      port map(D => un1_readmemoryaddrcounter_cry_2_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemoryaddrcounter_Z(29));
    
    \SPITransmitReg_RNO_0[29]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(21), Y => N_4_2);
    
    \ControllUnitState_RNO[0]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => ControllUnitState_ns_i_0_a2_0_1_Z(14), B => 
        N_4353, C => N_765, D => ControllUnitState_ns_i_0_0_Z(14), 
        Y => N_2554_i);
    
    \SPITransmitReg[31]\ : SLE
      port map(D => SPITransmitReg_13(31), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(31));
    
    \CurrentAddrReg[17]\ : SLE
      port map(D => un1_currentaddrreg_cry_17_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(17));
    
    \Stamp1ShadowReg2[16]\ : SLE
      port map(D => STAMP_0_data_frame(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(16));
    
    \StampFSMR1[1]\ : SLE
      port map(D => pageaddr_5_i_m4(1), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(1));
    
    \SPITransmitReg_RNO_0[22]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(14), Y => N_4_9);
    
    \mainProcess.PRDATA_8_0_iv_0[10]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(10), B => 
        PRDATA_8_0_iv_0_3(10), C => PRDATA_8_0_iv_0_6(10), Y => 
        PRDATA_8(10));
    
    \mainProcess.InternalData2Memory_27_0_iv[27]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_2(27), C => 
        Stamp1ShadowReg2_Z(27), D => 
        InternalData2Memory_27_0_iv_0(27), Y => 
        InternalData2Memory_27(27));
    
    \mainProcess.PRDATA_8_0_iv_0_3[11]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(11), B => 
        Stamp1ShadowReg2_Z(11), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(11));
    
    \mainProcess.PRDATA_8_0_iv_0_3[31]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(31), B => 
        Stamp1ShadowReg2_Z(31), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(31));
    
    \SPITransmitReg_RNO[30]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_1, B => InternalDataFromMem(30), C => 
        N_54, D => N_15_mux_0, Y => SPITransmitReg_13(30));
    
    \mainProcess.PRDATA_8_0_iv_0_2[18]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(18), 
        D => CurrentAddrReg_Z(18), Y => PRDATA_8_0_iv_0_2(18));
    
    un1_readmemoryaddrcounter_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemoryaddrcounter_Z(26), C
         => \GND\, D => \GND\, FCI => 
        un1_readmemoryaddrcounter_cry_4_Z, S => 
        un1_readmemoryaddrcounter_cry_5_S, Y => 
        un1_readmemoryaddrcounter_cry_5_Y, FCO => 
        un1_readmemoryaddrcounter_cry_5_Z);
    
    \memorycnt[4]\ : SLE
      port map(D => memorycnt_6(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => memorycnt_Z(4));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[7]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(7), C => 
        Stamp1ShadowReg2_Z(7), D => 
        InternalData2Memory_27_0_iv_0_1(7), Y => 
        InternalData2Memory_27(7));
    
    un1_currentaddrreg_cry_25 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(25), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_24_Z, S => 
        un1_currentaddrreg_cry_25_S, Y => 
        un1_currentaddrreg_cry_25_Y, FCO => 
        un1_currentaddrreg_cry_25_Z);
    
    InternalAddr2Memory_0_sqmuxa_i : CFG4
      generic map(INIT => x"FBBB")

      port map(A => APB3ReadMemoryLimitedState_RNI12J4_Y(5), B
         => N_138, C => InternalAddr2Memory_0_sqmuxa_2_i_a2_8_Z, 
        D => InternalAddr2Memory_0_sqmuxa_2_i_a2_7_Z, Y => 
        InternalAddr2Memory_0_sqmuxa_i_Z);
    
    \ReadMemoryState_ns_i_0_a3[3]\ : CFG4
      generic map(INIT => x"0301")

      port map(A => ReadMemoryState_Z(6), B => 
        ReadMemoryState_Z(5), C => ReadMemoryState_Z(4), D => 
        N_4274, Y => N_80);
    
    \mainProcess.InternalData2Memory_27_0_iv[30]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_2(30), C => 
        Stamp1ShadowReg2_Z(30), D => 
        InternalData2Memory_27_0_iv_0(30), Y => 
        InternalData2Memory_27(30));
    
    \ReadMemoryShadowReg[7]\ : SLE
      port map(D => InternalDataFromMem(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(7));
    
    \InternalAddr2Memory[1]\ : SLE
      port map(D => InternalAddr2Memory_34(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => InternalAddr2Memory_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => InternalAddr2Memory_Z(1));
    
    \APBState_ns_1_0_.m3_0_a2\ : CFG3
      generic map(INIT => x"02")

      port map(A => sb_sb_0_Memory_PSELx, B => N_1539_i, C => 
        sb_sb_0_STAMP_PWRITE, Y => APBState_ns(0));
    
    \readmemorylimitedcnt_RNI4GJ84[2]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => readmemorylimitedcnt_Z(2), B => 
        readmemorylimitedcnt_Z(7), C => m60_e_5, D => m60_e_4, Y
         => N_139_mux);
    
    \mainProcess.PRDATA_8_0_iv_0_a2_8[12]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => sb_sb_0_STAMP_PADDR(2), B => 
        sb_sb_0_STAMP_PADDR(4), C => sb_sb_0_STAMP_PADDR(6), D
         => sb_sb_0_STAMP_PADDR(5), Y => N_1030);
    
    \ControllUnitState_ns_0_0[5]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => ControllUnitState_Z(9), B => 
        ControllUnitState_Z(12), C => N_1045, D => N_712, Y => 
        ControllUnitState_ns(5));
    
    \CommandReg[28]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(28));
    
    un8_tempcounter_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => StampFSMPC_Z(4), C => \GND\, D
         => \GND\, FCI => un8_tempcounter_cry_3_Z, S => 
        un8_tempcounter_cry_4_S, Y => un8_tempcounter_cry_4_Y, 
        FCO => un8_tempcounter_cry_4_Z);
    
    \mainProcess.InternalAddr2Memory_34_18\ : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory_34_sm0, B => 
        InternalAddr2Memory_34_m0(2), C => N_143_mux, Y => 
        InternalAddr2Memory_34_18);
    
    \mainProcess.PRDATA_8_0_iv_0_3[26]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(26), B => 
        Stamp1ShadowReg2_Z(26), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(26));
    
    \InternalData2Memory[3]\ : SLE
      port map(D => InternalData2Memory_27(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(3));
    
    \SPITransmitReg[3]\ : SLE
      port map(D => SPITransmitReg_13(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(3));
    
    \StartAddrReg[6]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(6));
    
    \Stamp1ShadowReg1[11]\ : SLE
      port map(D => STAMP_0_data_frame(43), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(11));
    
    \readmemoryaddrcounter[27]\ : SLE
      port map(D => un1_readmemoryaddrcounter_cry_4_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemoryaddrcounter_Z(27));
    
    \StampFSMR1[0]\ : SLE
      port map(D => pageaddr_5_i_m4(0), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(0));
    
    \mainProcess.SPITransmitReg_13_0_iv_0_a2_2[30]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_4272_i, B => ReadMemoryState_Z(7), Y => 
        N_1034);
    
    \mainProcess.SPIaddr_15_iv_0[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => ConfigStatusReg_Z(0), B => N_4358, C => 
        SPIaddr_3_sqmuxa_1, Y => SPIaddr_15(0));
    
    \mainProcess.pageaddr_5_i_m4[28]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(28), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(28), Y => pageaddr_5_i_m4(28));
    
    \PRDATA[26]\ : SLE
      port map(D => PRDATA_8(26), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(26));
    
    \ControllUnitState_ns_0_0_o2[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => dataReady_0, B => ControllUnitState_Z(14), Y
         => N_4344);
    
    \un23_o2[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_4343_i, B => ControllUnitState_Z(4), Y => 
        N_1260);
    
    \mainProcess.InternalAddr2Memory_34_1[7]\ : CFG4
      generic map(INIT => x"0F44")

      port map(A => readmemoryaddrcounter_Z(24), B => 
        ReadMemoryState_Z(4), C => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), D => N_138, Y
         => InternalAddr2Memory_34_1(7));
    
    \SPITransmitReg_RNO_1[21]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(21), Y => N_15_mux_9);
    
    \mainProcess.PRDATA_8_0_iv_0_2[24]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(24), 
        D => CurrentAddrReg_Z(24), Y => PRDATA_8_0_iv_0_2(24));
    
    \ControllUnitState[6]\ : SLE
      port map(D => ControllUnitState_ns(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(6));
    
    \mainProcess.PRDATA_8_0_iv_0_0[20]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(20), D => SPIRecReg(20), Y => 
        PRDATA_8_0_iv_0_0(20));
    
    \mainProcess.PRDATA_8_0_iv_0[7]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(7), B => 
        PRDATA_8_0_iv_0_3(7), C => PRDATA_8_0_iv_0_6(7), Y => 
        PRDATA_8(7));
    
    \StartAddrReg[11]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(11));
    
    \APB3ReadMemoryLimitedState[0]\ : SLE
      port map(D => N_145_mux, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \GND\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => 
        APB3ReadMemoryLimitedState_Z(0));
    
    un1_readmemoryaddrcounter_s_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemoryaddrcounter_Z(23), C
         => \GND\, D => \GND\, FCI => 
        un1_readmemoryaddrcounter_cry_7_Z, S => 
        un1_readmemoryaddrcounter_s_8_S, Y => 
        un1_readmemoryaddrcounter_s_8_Y, FCO => 
        un1_readmemoryaddrcounter_s_8_FCO);
    
    \mainProcess.PRDATA_8_0_iv_0[26]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(26), B => 
        PRDATA_8_0_iv_0_3(26), C => PRDATA_8_0_iv_0_6(26), Y => 
        PRDATA_8(26));
    
    \ControllUnitState_ns_i_a5_i_o2[2]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_2624, B => ControllUnitState_Z(3), Y => 
        N_4349);
    
    \CurrentAddrReg[25]\ : SLE
      port map(D => un1_currentaddrreg_cry_25_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(25));
    
    ControllUnitState_tr25_0_a2_5 : CFG4
      generic map(INIT => x"0200")

      port map(A => tempcounter_Z(7), B => tempcounter_Z(3), C
         => tempcounter_Z(1), D => tempcounter_Z(0), Y => 
        ControllUnitState_tr25_0_a2_5_Z);
    
    \tempcounter[6]\ : SLE
      port map(D => N_4298_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_enabletimestampgen2_1_i, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tempcounter_Z(6));
    
    \StartAddrReg[20]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(20));
    
    \ControllUnitSubState_ns_0_a2_0[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => ControllUnitSubState_Z(0), B => 
        ControllUnitState_Z(3), Y => N_2648);
    
    \SPIState_RNO_2[4]\ : CFG3
      generic map(INIT => x"10")

      port map(A => SPIState_Z(0), B => SPIState_Z(2), C => m46_0, 
        Y => m46_1_1_0_1);
    
    \mainProcess.InternalData2Memory_27_0_iv_0[11]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(11), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0(11));
    
    \mainProcess.InternalData2Memory_27_0_iv_1[21]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0(21), C => pageaddr(29), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_1(21));
    
    \SPITransmitReg_RNO_0[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(3), Y => N_4_20);
    
    \ControllUnitState_ns_0_0_a2[5]\ : CFG4
      generic map(INIT => x"8400")

      port map(A => ControllUnitSubState_Z(1), B => dataReady_0, 
        C => ControllUnitSubState_Z(0), D => 
        ControllUnitState_Z(3), Y => N_712);
    
    \Stamp1ShadowReg2[20]\ : SLE
      port map(D => STAMP_0_data_frame(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(20));
    
    \ControllUnitState_ns_i_a5_i[2]\ : CFG4
      generic map(INIT => x"FF10")

      port map(A => N_4339, B => N_4349, C => dataReady_0, D => 
        ControllUnitState_Z(10), Y => N_161);
    
    \mainProcess.PRDATA_8_0_iv_0_0[22]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(22), D => SPIRecReg(22), Y => 
        PRDATA_8_0_iv_0_0(22));
    
    \ControllUnitSubState_RNI80EH[0]\ : CFG4
      generic map(INIT => x"0B00")

      port map(A => ControllUnitSubState_Z(0), B => 
        ControllUnitState_Z(2), C => ConfigStatusReg_24_sn_N_5, D
         => GPIO_6_M2F_c, Y => un1_enabletimestampgen2_1_i);
    
    un1_APBState_1_1_0_a2_0 : CFG3
      generic map(INIT => x"04")

      port map(A => sb_sb_0_STAMP_PADDR(6), B => N_1028, C => 
        sb_sb_0_STAMP_PADDR(2), Y => N_4547);
    
    \SPIState_RNO_0[0]\ : CFG2
      generic map(INIT => x"7")

      port map(A => N_21_0, B => m33_e_0, Y => N_154_mux_i_1_0);
    
    \mainProcess.PRDATA_8_0_iv_0[29]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(29), B => 
        PRDATA_8_0_iv_0_3(29), C => PRDATA_8_0_iv_0_6(29), Y => 
        PRDATA_8(29));
    
    \InternalData2Memory[18]\ : SLE
      port map(D => InternalData2Memory_27(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(18));
    
    \CommandReg[18]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(18));
    
    \ReadMemoryState_RNO_0[8]\ : CFG4
      generic map(INIT => x"035F")

      port map(A => N_4274, B => N_68, C => ReadMemoryState_Z(6), 
        D => N_62, Y => N_2471_i_1);
    
    \mainProcess.PRDATA_8_0_iv_0_0[23]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(23), D => SPIRecReg(23), Y => 
        PRDATA_8_0_iv_0_0(23));
    
    \mainProcess.PRDATA_8_0_iv_0_2[9]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(9), 
        D => CurrentAddrReg_Z(9), Y => PRDATA_8_0_iv_0_2(9));
    
    \readmemorycounter_RNO[3]\ : CFG4
      generic map(INIT => x"3120")

      port map(A => un1_enableSPI_1_sqmuxa_1_i, B => N_95, C => 
        N_4274, D => N_1508_i, Y => N_4262_i);
    
    MemoryPageSize_1_sqmuxa_0_o4_0 : CFG4
      generic map(INIT => x"DFFF")

      port map(A => APBState_Z(1), B => sb_sb_0_STAMP_PADDR(3), C
         => sb_sb_0_STAMP_PADDR(2), D => sb_sb_0_STAMP_PADDR(6), 
        Y => MemoryPageSize_1_sqmuxa_0_o4_0_Z);
    
    \StampFSMR1[13]\ : SLE
      port map(D => pageaddr_5_i_m4(13), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(13));
    
    \mainProcess.PRDATA_8_0_iv_0_1[25]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ConfigStatusReg_Z(25), B => CommandReg_Z(25), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(25));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[22]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(22), C => pageaddr(30), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(22));
    
    \mainProcess.InternalData2Memory_27_0_iv_3[25]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(25), B => 
        TimeStampValue(25), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_3(25));
    
    Command_1_sqmuxa_0_a2_0 : CFG3
      generic map(INIT => x"40")

      port map(A => sb_sb_0_STAMP_PADDR(2), B => 
        sb_sb_0_STAMP_PADDR(6), C => sb_sb_0_STAMP_PADDR(3), Y
         => N_1025);
    
    \SPITransmitReg_RNO_1[15]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(15), Y => N_15_mux_15);
    
    \mainProcess.PRDATA_8_0_iv_0_6[6]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(6), C => 
        PRDATA_8_0_iv_0_1(6), D => PRDATA_8_0_iv_0_0(6), Y => 
        PRDATA_8_0_iv_0_6(6));
    
    \ControllUnitSubState_ns_0_0_a2_1_2[0]\ : CFG3
      generic map(INIT => x"40")

      port map(A => ControllUnitState_Z(2), B => N_1041, C => 
        ControllUnitSubState_Z(0), Y => 
        ControllUnitSubState_ns_0_0_a2_1_Z(0));
    
    \SPITransmitReg_RNO[29]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_2, B => InternalDataFromMem(29), C => 
        N_54, D => N_15_mux_1, Y => SPITransmitReg_13(29));
    
    \mainProcess.pageaddr_5_i_m4[17]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(17), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(17), Y => N_4371);
    
    un1_enabletimestampgen2_5_8 : CFG4
      generic map(INIT => x"FFE0")

      port map(A => ControllUnitState_Z(5), B => 
        ControllUnitState_Z(6), C => N_4343_i, D => 
        un1_enabletimestampgen2_5_6_Z, Y => 
        un1_enabletimestampgen2_5_8_Z);
    
    \InternalAddr2Memory[0]\ : SLE
      port map(D => InternalAddr2Memory_34(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => InternalAddr2Memory_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => InternalAddr2Memory_Z(0));
    
    \SPIState_RNO_3[4]\ : CFG4
      generic map(INIT => x"40C0")

      port map(A => SPIState_Z(2), B => m46_0, C => m33_e_0, D
         => counter9, Y => m46_1_1_tz);
    
    \ReadMemoryState[0]\ : SLE
      port map(D => ReadMemoryState_ns_i_i_Z(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \GND\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ReadMemoryState_Z(0));
    
    un1_currentaddrreg_cry_2 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(2), B => pageaddr(2), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_1_Z, S
         => un1_currentaddrreg_cry_2_S, Y => 
        un1_currentaddrreg_cry_2_Y, FCO => 
        un1_currentaddrreg_cry_2_Z);
    
    \ControllUnitSubState_ns_i_a7_0_2[1]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => ControllUnitState_Z(7), B => 
        ControllUnitState_Z(8), C => ControllUnitSubState_Z(0), D
         => ControllUnitState_Z(9), Y => 
        ControllUnitSubState_ns_i_a7_0_2_Z(1));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[3]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(3), B => TimeStampValue(3), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(3));
    
    \mainProcess.InternalAddr2Memory_34_2\ : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory_34_sm0, B => 
        InternalAddr2Memory_34_m0(5), C => N_143_mux, Y => 
        InternalAddr2Memory_34_2);
    
    InternalAddr2Memory_0_sqmuxa_2_i_a2_1 : CFG4
      generic map(INIT => x"0001")

      port map(A => ControllUnitState_Z(12), B => 
        ControllUnitState_Z(0), C => ControllUnitState_Z(14), D
         => ControllUnitState_Z(1), Y => 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_1_Z);
    
    \StampFSMR1[17]\ : SLE
      port map(D => N_4371, CLK => sb_sb_0_FIC_0_CLK, EN => 
        ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        pageaddr(17));
    
    \Stamp1ShadowReg1[5]\ : SLE
      port map(D => STAMP_0_data_frame(37), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(5));
    
    \mainProcess.PRDATA_8_0_iv_0_2[11]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(11), 
        D => CurrentAddrReg_Z(11), Y => PRDATA_8_0_iv_0_2(11));
    
    \StartAddrReg[19]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(19));
    
    \mainProcess.SPIaddr_15_iv_0_m2[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => ConfigStatusReg_Z(31), B => 
        SPIaddr_0_sqmuxa_3, C => N_155_mux_i, Y => N_4358);
    
    \mainProcess.pageaddr_5_i_m4[13]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(13), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(13), Y => pageaddr_5_i_m4(13));
    
    un1_enabletimestampgen2_5_2 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => ControllUnitState_Z(14), B => 
        ControllUnitState_Z(2), C => ControllUnitState_Z(13), D
         => ControllUnitState_Z(12), Y => 
        un1_enabletimestampgen2_5_2_Z);
    
    \InternalAddr2Memory[5]\ : SLE
      port map(D => InternalAddr2Memory_34(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => InternalAddr2Memory_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => InternalAddr2Memory_Z(5));
    
    un1_currentaddrreg_cry_8 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(8), B => pageaddr(8), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_7_Z, S
         => un1_currentaddrreg_cry_8_S, Y => 
        un1_currentaddrreg_cry_8_Y, FCO => 
        un1_currentaddrreg_cry_8_Z);
    
    \StampFSMR1[24]\ : SLE
      port map(D => pageaddr_5_i_m4(24), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(24));
    
    \SPITransmitReg[7]\ : SLE
      port map(D => SPITransmitReg_13(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(7));
    
    \SPITransmitReg_RNO[23]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_8, B => InternalDataFromMem(23), C => 
        N_54, D => N_15_mux_7, Y => SPITransmitReg_13(23));
    
    \mainProcess.PRDATA_8_0_iv_0_3[28]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(28), B => 
        Stamp1ShadowReg2_Z(28), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(28));
    
    \CommandReg[20]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(20));
    
    \mainProcess.PRDATA_8_0_iv_0_3[0]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(0), B => 
        Stamp1ShadowReg2_Z(0), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(0));
    
    InternalData2Memory_3_sqmuxa : CFG2
      generic map(INIT => x"1")

      port map(A => N_1232_i, B => ReadMemoryState_Z(4), Y => 
        InternalData2Memory_3_sqmuxa_Z);
    
    \mainProcess.PRDATA_8_0_iv_0_1[16]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(8), B => CommandReg_Z(16), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(16));
    
    enableSPI_0_sqmuxa_2_0_a2 : CFG4
      generic map(INIT => x"001D")

      port map(A => SPIState_Z(3), B => SPIState_Z(2), C => N_144, 
        D => N_62, Y => enableSPI_0_sqmuxa_2);
    
    \mainProcess.PRDATA_8_0_iv_0_6[2]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(2), C => 
        PRDATA_8_0_iv_0_1(2), D => PRDATA_8_0_iv_0_0(2), Y => 
        PRDATA_8_0_iv_0_6(2));
    
    \SPITransmitReg[0]\ : SLE
      port map(D => SPITransmitReg_13(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(0));
    
    \readmemorylimitedcnt_RNICOMS1[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => readmemorylimitedcnt_Z(5), B => 
        readmemorylimitedcnt_Z(4), C => readmemorylimitedcnt_Z(3), 
        D => readmemorylimitedcnt_Z(0), Y => m60_e_5);
    
    \mainProcess.PRDATA_8_0_iv_0_0[9]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(9), D => SPIRecReg(9), Y => 
        PRDATA_8_0_iv_0_0(9));
    
    \ReadMemoryShadowReg[23]\ : SLE
      port map(D => InternalDataFromMem(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(23));
    
    \ControllUnitSubState_ns_i_1[1]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ControllUnitSubState_Z(0), B => 
        ControllUnitSubState_ns_i_0_Z(1), C => dataReady_0, D => 
        ControllUnitState_Z(3), Y => 
        ControllUnitSubState_ns_i_1_Z(1));
    
    \StartAddrReg[18]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(18));
    
    \SPIState_RNO_1[4]\ : CFG3
      generic map(INIT => x"2E")

      port map(A => SPIState_Z(0), B => SPIState_Z(2), C => 
        counter9, Y => m46_1_1);
    
    \mainProcess.PRDATA_8_0_iv_0_0[19]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(19), D => SPIRecReg(19), Y => 
        PRDATA_8_0_iv_0_0(19));
    
    \mainProcess.readmemorylimitedcnt_5_RNO[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemorylimitedcnt_Z(8), C => 
        \GND\, D => \GND\, FCI => un1_readmemorylimitedcnt_cry_7, 
        S => readmemorylimitedcnt_5_RNO_S(8), Y => 
        readmemorylimitedcnt_5_RNO_Y(8), FCO => 
        readmemorylimitedcnt_5_RNO_FCO(8));
    
    \mainProcess.PRDATA_8_0_iv_0[18]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(18), B => 
        PRDATA_8_0_iv_0_3(18), C => PRDATA_8_0_iv_0_6(18), Y => 
        PRDATA_8(18));
    
    \CommandReg[30]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(30));
    
    \SPIState[1]\ : SLE
      port map(D => SPIState_ns(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => SPIState_Z(1));
    
    SPI : spi_master_2_32
      port map(SPITransmitReg(31) => SPITransmitReg_Z(31), 
        SPITransmitReg(30) => SPITransmitReg_Z(30), 
        SPITransmitReg(29) => SPITransmitReg_Z(29), 
        SPITransmitReg(28) => SPITransmitReg_Z(28), 
        SPITransmitReg(27) => SPITransmitReg_Z(27), 
        SPITransmitReg(26) => SPITransmitReg_Z(26), 
        SPITransmitReg(25) => SPITransmitReg_Z(25), 
        SPITransmitReg(24) => SPITransmitReg_Z(24), 
        SPITransmitReg(23) => SPITransmitReg_Z(23), 
        SPITransmitReg(22) => SPITransmitReg_Z(22), 
        SPITransmitReg(21) => SPITransmitReg_Z(21), 
        SPITransmitReg(20) => SPITransmitReg_Z(20), 
        SPITransmitReg(19) => SPITransmitReg_Z(19), 
        SPITransmitReg(18) => SPITransmitReg_Z(18), 
        SPITransmitReg(17) => SPITransmitReg_Z(17), 
        SPITransmitReg(16) => SPITransmitReg_Z(16), 
        SPITransmitReg(15) => SPITransmitReg_Z(15), 
        SPITransmitReg(14) => SPITransmitReg_Z(14), 
        SPITransmitReg(13) => SPITransmitReg_Z(13), 
        SPITransmitReg(12) => SPITransmitReg_Z(12), 
        SPITransmitReg(11) => SPITransmitReg_Z(11), 
        SPITransmitReg(10) => SPITransmitReg_Z(10), 
        SPITransmitReg(9) => SPITransmitReg_Z(9), 
        SPITransmitReg(8) => SPITransmitReg_Z(8), 
        SPITransmitReg(7) => SPITransmitReg_Z(7), 
        SPITransmitReg(6) => SPITransmitReg_Z(6), 
        SPITransmitReg(5) => SPITransmitReg_Z(5), 
        SPITransmitReg(4) => SPITransmitReg_Z(4), 
        SPITransmitReg(3) => SPITransmitReg_Z(3), 
        SPITransmitReg(2) => SPITransmitReg_Z(2), 
        SPITransmitReg(1) => SPITransmitReg_Z(1), 
        SPITransmitReg(0) => SPITransmitReg_Z(0), SPIaddr_0 => 
        SPIaddr_Z(0), SPIRecReg(31) => SPIRecReg(31), 
        SPIRecReg(30) => SPIRecReg(30), SPIRecReg(29) => 
        SPIRecReg(29), SPIRecReg(28) => SPIRecReg(28), 
        SPIRecReg(27) => SPIRecReg(27), SPIRecReg(26) => 
        SPIRecReg(26), SPIRecReg(25) => SPIRecReg(25), 
        SPIRecReg(24) => SPIRecReg(24), SPIRecReg(23) => 
        SPIRecReg(23), SPIRecReg(22) => SPIRecReg(22), 
        SPIRecReg(21) => SPIRecReg(21), SPIRecReg(20) => 
        SPIRecReg(20), SPIRecReg(19) => SPIRecReg(19), 
        SPIRecReg(18) => SPIRecReg(18), SPIRecReg(17) => 
        SPIRecReg(17), SPIRecReg(16) => SPIRecReg(16), 
        SPIRecReg(15) => SPIRecReg(15), SPIRecReg(14) => 
        SPIRecReg(14), SPIRecReg(13) => SPIRecReg(13), 
        SPIRecReg(12) => SPIRecReg(12), SPIRecReg(11) => 
        SPIRecReg(11), SPIRecReg(10) => SPIRecReg(10), 
        SPIRecReg(9) => SPIRecReg(9), SPIRecReg(8) => 
        SPIRecReg(8), SPIRecReg(7) => SPIRecReg(7), SPIRecReg(6)
         => SPIRecReg(6), SPIRecReg(5) => SPIRecReg(5), 
        SPIRecReg(4) => SPIRecReg(4), SPIRecReg(3) => 
        SPIRecReg(3), SPIRecReg(2) => SPIRecReg(2), SPIRecReg(1)
         => SPIRecReg(1), SPIRecReg(0) => SPIRecReg(0), enable
         => enable, InternalBusy => InternalBusy, mosi_cl_1z => 
        mosi_cl, mosi_1_1z => mosi_1, resetn => resetn, SCLK_c
         => SCLK_c, MISO_c => MISO_c, nCS2_c => nCS2_c, 
        resetn_arst => resetn_arst, nCS1_c => nCS1_c, 
        sb_sb_0_FIC_0_CLK => sb_sb_0_FIC_0_CLK);
    
    PREADY : SLE
      port map(D => N_1539_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        resetn, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => sb_sb_0_Memory_PREADY);
    
    \readmemoryaddrcounter[28]\ : SLE
      port map(D => un1_readmemoryaddrcounter_cry_3_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemoryaddrcounter_Z(28));
    
    \PRDATA[7]\ : SLE
      port map(D => PRDATA_8(7), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(7));
    
    \Stamp1ShadowReg1[14]\ : SLE
      port map(D => STAMP_0_data_frame(46), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(14));
    
    \SPITransmitReg_RNO_1[19]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(19), Y => N_15_mux_11);
    
    \SPITransmitReg[24]\ : SLE
      port map(D => SPITransmitReg_13(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(24));
    
    \SPITransmitReg[22]\ : SLE
      port map(D => SPITransmitReg_13(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(22));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_a2_0[28]\ : CFG3
      generic map(INIT => x"40")

      port map(A => ReadMemoryState_Z(4), B => pageaddr(4), C => 
        ControllUnitState_Z(10), Y => N_4535);
    
    InternalData2Memory_4_sqmuxa : CFG3
      generic map(INIT => x"04")

      port map(A => N_1255_i, B => ControllUnitState_Z(9), C => 
        ReadMemoryState_Z(4), Y => InternalData2Memory_4_sqmuxa_Z);
    
    \mainProcess.InternalData2Memory_27_0_iv_1[11]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0(11), C => pageaddr(19), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_1(11));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[16]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(16), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(16));
    
    StartAddrReg_0_sqmuxa_0_a2 : CFG3
      generic map(INIT => x"20")

      port map(A => N_1186, B => sb_sb_0_STAMP_PADDR(6), C => 
        N_1029, Y => StartAddrReg_0_sqmuxa);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[12]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(12), C => pageaddr(20), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(12));
    
    un8_tempcounter_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => StampFSMPC_Z(5), C => \GND\, D
         => \GND\, FCI => un8_tempcounter_cry_4_Z, S => 
        un8_tempcounter_cry_5_S, Y => un8_tempcounter_cry_5_Y, 
        FCO => un8_tempcounter_cry_5_Z);
    
    \InternalData2Memory[7]\ : SLE
      port map(D => InternalData2Memory_27(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(7));
    
    \SPITransmitReg_RNO_1[12]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(12), Y => N_15_mux_18);
    
    \Stamp1ShadowReg2[11]\ : SLE
      port map(D => STAMP_0_data_frame(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(11));
    
    \Command_RNO[6]\ : CFG2
      generic map(INIT => x"2")

      port map(A => sb_sb_0_STAMP_PWDATA(30), B => 
        SPIState_RNI27U44_Z(1), Y => N_168_i);
    
    \mainProcess.ConfigStatusReg_26_0_m2_1[30]\ : CFG3
      generic map(INIT => x"53")

      port map(A => ConfigStatusReg_Z(30), B => N_1316_i, C => 
        N_4354, Y => ConfigStatusReg_26_0_m2_1(30));
    
    \Stamp1ShadowReg1[27]\ : SLE
      port map(D => STAMP_0_data_frame(59), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(27));
    
    \ConfigStatusReg_RNO_1[4]\ : CFG3
      generic map(INIT => x"31")

      port map(A => N_81, B => ReadMemoryState_Z(3), C => 
        APB3ReadMemoryLimitedState_Z(1), Y => d_N_5_mux);
    
    \StampFSMPC_6_0_a2[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => un8_tempcounter_cry_5_S, B => 
        ControllUnitState_Z(11), Y => StampFSMPC_6(5));
    
    \mainProcess.PRDATA_8_0_iv_0_6[27]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(27), C => 
        PRDATA_8_0_iv_0_1(27), D => PRDATA_8_0_iv_0_0(27), Y => 
        PRDATA_8_0_iv_0_6(27));
    
    un1_enabletimestampgen2_7_0_0 : CFG4
      generic map(INIT => x"01FF")

      port map(A => ControllUnitState_Z(9), B => 
        ControllUnitSubState_Z(1), C => ControllUnitState_Z(11), 
        D => GPIO_6_M2F_c, Y => un1_enabletimestampgen2_7_0_0_Z);
    
    \InternalAddr2Memory[8]\ : SLE
      port map(D => InternalAddr2Memory_34(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => InternalAddr2Memory_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => InternalAddr2Memory_Z(8));
    
    \SPIState_RNITHKL1[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => counter9, B => SPIState_Z(2), Y => 
        SPIState_ns(3));
    
    \PRDATA[14]\ : SLE
      port map(D => PRDATA_8(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(14));
    
    \StartAddrReg[1]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(1));
    
    \mainProcess.InternalData2Memory_27_0_iv_2[24]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(24), B => 
        TimeStampValue(24), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_2(24));
    
    \mainProcess.PRDATA_8_0_iv_0_6[19]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(19), C => 
        PRDATA_8_0_iv_0_1(19), D => PRDATA_8_0_iv_0_0(19), Y => 
        PRDATA_8_0_iv_0_6(19));
    
    InternalAddr2Memory_0_sqmuxa_2_i_a2_7 : CFG4
      generic map(INIT => x"10F0")

      port map(A => ControllUnitState_Z(5), B => 
        ControllUnitState_Z(7), C => GPIO_6_M2F_c, D => N_4343_i, 
        Y => InternalAddr2Memory_0_sqmuxa_2_i_a2_7_Z);
    
    \ControllUnitState_ns_i_0_a2_0_1[14]\ : CFG2
      generic map(INIT => x"1")

      port map(A => ControllUnitState_Z(14), B => 
        ControllUnitState_Z(0), Y => N_765_1);
    
    \CommandReg[10]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(10));
    
    \SPITransmitReg_RNO_0[23]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(15), Y => N_4_8);
    
    \mainProcess.PRDATA_8_0_iv_0_0[24]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(24), D => SPIRecReg(24), Y => 
        PRDATA_8_0_iv_0_0(24));
    
    \StampFSMR1[6]\ : SLE
      port map(D => pageaddr_5_i_m4(6), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(6));
    
    \StampFSMR1[2]\ : SLE
      port map(D => pageaddr_5_i_m4(2), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(2));
    
    \mainProcess.SPITransmitReg_13_0_iv_0[5]\ : CFG4
      generic map(INIT => x"A808")

      port map(A => N_4270, B => InternalDataFromMem(5), C => 
        SPIState_1_sqmuxa, D => sb_sb_0_STAMP_PWDATA(5), Y => 
        SPITransmitReg_13(5));
    
    \mainProcess.InternalAddr2Memory_34[7]\ : CFG4
      generic map(INIT => x"DCDD")

      port map(A => InternalAddr2Memory_34_1(7), B => 
        InternalAddr2Memory_34_10, C => readmemorylimitedcnt_Z(7), 
        D => N_138, Y => InternalAddr2Memory_34(7));
    
    \SPITransmitReg_RNO_0[30]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(22), Y => N_4_1);
    
    \mainProcess.tempcounter_7_iv_i[0]\ : CFG3
      generic map(INIT => x"0B")

      port map(A => N_1261_i, B => StampFSMPC_Z(0), C => 
        ControllUnitState_Z(1), Y => tempcounter_7_iv_i(0));
    
    \InternalData2Memory[6]\ : SLE
      port map(D => InternalData2Memory_27(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(6));
    
    \InternalAddr2Memory[7]\ : SLE
      port map(D => InternalAddr2Memory_34(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => InternalAddr2Memory_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => InternalAddr2Memory_Z(7));
    
    \Stamp1ShadowReg1[23]\ : SLE
      port map(D => STAMP_0_data_frame(55), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(23));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[1]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(1), C => 
        Stamp1ShadowReg2_Z(1), D => 
        InternalData2Memory_27_0_iv_0_1(1), Y => 
        InternalData2Memory_27(1));
    
    \mainProcess.PRDATA_8_0_iv_0[9]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(9), B => 
        PRDATA_8_0_iv_0_3(9), C => PRDATA_8_0_iv_0_6(9), Y => 
        PRDATA_8(9));
    
    \ControllUnitState[11]\ : SLE
      port map(D => ControllUnitState_Z(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(11));
    
    \CurrentAddrReg[1]\ : SLE
      port map(D => un1_currentaddrreg_cry_1_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(1));
    
    \ReadMemoryState_ns_i_i[8]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => ReadMemoryState_Z(1), B => 
        ReadMemoryState_Z(0), C => N_2496, Y => 
        ReadMemoryState_ns_i_i_Z(8));
    
    WriteEnable_0_sqmuxa_i : CFG4
      generic map(INIT => x"FFF1")

      port map(A => N_1302, B => un1_enabletimestampgen2_7_0_0_Z, 
        C => ReadMemoryState_Z(5), D => ReadMemoryState_Z(4), Y
         => WriteEnable_0_sqmuxa_i_Z);
    
    un1_APBState_1_2_0 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => sb_sb_0_STAMP_PADDR(9), B => 
        sb_sb_0_STAMP_PADDR(8), C => sb_sb_0_STAMP_PADDR(7), D
         => sb_sb_0_STAMP_PADDR(10), Y => un1_APBState_1_2_0_Z);
    
    \mainProcess.InternalAddr2Memory_34_6\ : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory_34_sm0, B => 
        InternalAddr2Memory_34_m0(4), C => N_143_mux, Y => 
        InternalAddr2Memory_34_6);
    
    \ControllUnitState_ns_0_0[7]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ControllUnitState_Z(8), B => 
        ControllUnitState_Z(7), C => N_4339, D => N_1045, Y => 
        ControllUnitState_ns(7));
    
    \ReadMemoryShadowReg[4]\ : SLE
      port map(D => InternalDataFromMem(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(4));
    
    \InternalData2Memory[30]\ : SLE
      port map(D => InternalData2Memory_27(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(30));
    
    \mainProcess.PRDATA_8_0_iv_0[4]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(4), B => 
        PRDATA_8_0_iv_0_3(4), C => PRDATA_8_0_iv_0_6(4), Y => 
        PRDATA_8(4));
    
    \mainProcess.PRDATA_8_0_iv_0_0[0]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(0), D => SPIRecReg(0), Y => 
        PRDATA_8_0_iv_0_0(0));
    
    \ReadMemoryState[3]\ : SLE
      port map(D => ReadMemoryState_ns(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ReadMemoryState_Z(3));
    
    InternalData2Memory_0_sqmuxa_6_i : CFG4
      generic map(INIT => x"F0F4")

      port map(A => un1_enabletimestampgen2_5_7_Z, B => 
        GPIO_6_M2F_c, C => ReadMemoryState_Z(4), D => 
        un1_enabletimestampgen2_5_8_Z, Y => 
        InternalData2Memory_0_sqmuxa_6_i_Z);
    
    \SPITransmitReg[20]\ : SLE
      port map(D => SPITransmitReg_13(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(20));
    
    \ControllUnitState_ns_0_0[12]\ : CFG4
      generic map(INIT => x"F2F0")

      port map(A => ControllUnitState_Z(2), B => 
        ConfigStatusReg_Z(2), C => N_734, D => N_4353, Y => 
        ControllUnitState_ns(12));
    
    \memorycnt[6]\ : SLE
      port map(D => memorycnt_6(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => memorycnt_Z(6));
    
    \SPITransmitReg_RNO_0[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(0), Y => N_4_23);
    
    \mainProcess.memorycnt_6_cry_0_0\ : ARI1
      generic map(INIT => x"5EDEE")

      port map(A => ControllUnitState_Z(3), B => memorycnt_Z(1), 
        C => ControllUnitState_RNI2VHT_Z(14), D => N_1255_i, FCI
         => \GND\, S => memorycnt_6_cry_0_0_S, Y => 
        memorycnt_6_cry_0_0_Y, FCO => memorycnt_6_cry_0);
    
    \StartAddrReg[3]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(3));
    
    \SPITransmitReg[13]\ : SLE
      port map(D => SPITransmitReg_13(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(13));
    
    \mainProcess.PRDATA_8_0_iv_0_1[9]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize(1), B => CommandReg_Z(9), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(9));
    
    \mainProcess.PRDATA_8_0_iv_0[1]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(1), B => 
        PRDATA_8_0_iv_0_3(1), C => PRDATA_8_0_iv_0_6(1), Y => 
        PRDATA_8(1));
    
    \Stamp1ShadowReg2[31]\ : SLE
      port map(D => STAMP_0_data_frame(31), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(31));
    
    \InternalData2Memory[17]\ : SLE
      port map(D => InternalData2Memory_27(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(17));
    
    \SPITransmitReg_RNO_0[4]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(4), Y => N_13_mux);
    
    \mainProcess.readmemorylimitedcnt_5[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => readmemorylimitedcnt_RNITM0U3_S(7), B => 
        APB3ReadMemoryLimitedState_Z(1), Y => 
        readmemorylimitedcnt_5(7));
    
    \mainProcess.PRDATA_8_0_iv_0[0]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(0), B => 
        PRDATA_8_0_iv_0_3(0), C => PRDATA_8_0_iv_0_6(0), Y => 
        PRDATA_8(0));
    
    \ControllUnitSubState[0]\ : SLE
      port map(D => ControllUnitSubState_ns(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitSubState_Z(0));
    
    \PRDATA[27]\ : SLE
      port map(D => PRDATA_8(27), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(27));
    
    \mainProcess.PRDATA_8_0_iv_0_1[8]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize(0), B => CommandReg_Z(8), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(8));
    
    \ReadMemoryShadowReg[16]\ : SLE
      port map(D => InternalDataFromMem(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(16));
    
    \mainProcess.PRDATA_8_0_iv_0_3[21]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(21), B => 
        Stamp1ShadowReg2_Z(21), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(21));
    
    \mainProcess.PRDATA_8_0_iv_0_2[31]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(31), 
        D => CurrentAddrReg_Z(31), Y => PRDATA_8_0_iv_0_2(31));
    
    ConfigStatusReg_2_sqmuxa_i_a3_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => ControllUnitState_Z(12), B => 
        ControllUnitState_Z(13), Y => N_1316_i);
    
    \mainProcess.PRDATA_8_0_iv_0_1[20]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(12), B => CommandReg_Z(20), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(20));
    
    \SPIState_RNI27U44[1]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => N_2496_i, B => N_71, C => SPIState_Z(1), Y
         => SPIState_RNI27U44_Z(1));
    
    \mainProcess.PRDATA_8_0_iv_0_2[7]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(7), 
        D => CurrentAddrReg_Z(7), Y => PRDATA_8_0_iv_0_2(7));
    
    \MemoryPageSize[12]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(12));
    
    \mainProcess.PRDATA_8_0_iv_0_2[5]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(5), 
        D => CurrentAddrReg_Z(5), Y => PRDATA_8_0_iv_0_2(5));
    
    un8_tempcounter_s_1_835 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => StampFSMPC_Z(0), C => \GND\, D
         => \GND\, FCI => \VCC\, S => un8_tempcounter_s_1_835_S, 
        Y => un8_tempcounter_s_1_835_Y, FCO => 
        un8_tempcounter_s_1_835_FCO);
    
    \mainProcess.PRDATA_8_0_iv_0_1[18]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(10), B => CommandReg_Z(18), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(18));
    
    \Command[2]\ : SLE
      port map(D => N_176_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        Command_1_sqmuxa_1_i_Z, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        Command_Z(2));
    
    un1_currentaddrreg_cry_21 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(21), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_20_Z, S => 
        un1_currentaddrreg_cry_21_S, Y => 
        un1_currentaddrreg_cry_21_Y, FCO => 
        un1_currentaddrreg_cry_21_Z);
    
    \PRDATA[28]\ : SLE
      port map(D => PRDATA_8(28), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(28));
    
    un8_tempcounter_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => StampFSMPC_Z(1), C => \GND\, D
         => \GND\, FCI => un8_tempcounter_s_1_835_FCO, S => 
        un8_tempcounter_cry_1_S, Y => un8_tempcounter_cry_1_Y, 
        FCO => un8_tempcounter_cry_1_Z);
    
    un1_currentaddrreg_cry_5 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(5), B => pageaddr(5), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_4_Z, S
         => un1_currentaddrreg_cry_5_S, Y => 
        un1_currentaddrreg_cry_5_Y, FCO => 
        un1_currentaddrreg_cry_5_Z);
    
    \StampFSMR1[30]\ : SLE
      port map(D => pageaddr_5_i_m4(30), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(30));
    
    \Stamp1ShadowReg1[26]\ : SLE
      port map(D => STAMP_0_data_frame(58), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(26));
    
    \CommandReg[24]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(24));
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    \SPITransmitReg_RNO[31]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_0, B => InternalDataFromMem(31), C => 
        N_54, D => N_15_mux, Y => SPITransmitReg_13(31));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[0]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(0), C => pageaddr(8), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(0));
    
    \ConfigStatusReg[8]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize(0));
    
    \Stamp1ShadowReg1[0]\ : SLE
      port map(D => STAMP_0_data_frame(32), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(0));
    
    \readmemorylimitedcnt[1]\ : SLE
      port map(D => readmemorylimitedcnt_5(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \GND\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorylimitedcnt_Z(1));
    
    \mainProcess.pageaddr_5_i_m4[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(4), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(4), Y => pageaddr_5_i_m4(4));
    
    \Command_RNO[2]\ : CFG2
      generic map(INIT => x"2")

      port map(A => sb_sb_0_STAMP_PWDATA(26), B => 
        SPIState_RNI27U44_Z(1), Y => N_176_i);
    
    \StampFSMR1[23]\ : SLE
      port map(D => pageaddr_5_i_m4(23), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(23));
    
    \un23_a3_0_0[1]\ : CFG4
      generic map(INIT => x"1110")

      port map(A => ControllUnitState_Z(6), B => 
        ControllUnitState_Z(5), C => ControllUnitSubState_Z(0), D
         => ControllUnitSubState_Z(1), Y => un23_a3_0(1));
    
    \SPITransmitReg_RNO[9]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_22, B => InternalDataFromMem(9), C => 
        N_54, D => N_15_mux_21, Y => SPITransmitReg_13(9));
    
    \InternalData2Memory[20]\ : SLE
      port map(D => InternalData2Memory_27(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(20));
    
    Command_1_sqmuxa_1_i_RNO_1 : CFG4
      generic map(INIT => x"0002")

      port map(A => APBState_Z(1), B => sb_sb_0_STAMP_PADDR(1), C
         => sb_sb_0_STAMP_PADDR(0), D => sb_sb_0_STAMP_PADDR(11), 
        Y => m73_m2_e_0_0);
    
    Command_1_sqmuxa_1_i_RNO : CFG3
      generic map(INIT => x"10")

      port map(A => sb_sb_0_STAMP_PADDR(9), B => 
        sb_sb_0_STAMP_PADDR(8), C => m73_m2_e_1, Y => m73_m2_e_2);
    
    un1_currentaddrreg_cry_15 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize(15), B => pageaddr(15), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_14_Z, S
         => un1_currentaddrreg_cry_15_S, Y => 
        un1_currentaddrreg_cry_15_Y, FCO => 
        un1_currentaddrreg_cry_15_Z);
    
    \tempcounter_RNO[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_1261_i, B => un8_tempcounter_cry_5_S, Y => 
        N_4297_i);
    
    \mainProcess.PRDATA_8_0_iv_0_3[9]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(9), B => 
        Stamp1ShadowReg2_Z(9), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(9));
    
    \mainProcess.PRDATA_8_0_iv_0_1[22]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize(14), B => CommandReg_Z(22), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(22));
    
    getTime : SLE
      port map(D => getTime_3, CLK => sb_sb_0_FIC_0_CLK, EN => 
        GPIO_6_M2F_c, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => getTime_Z);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[7]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(7), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(7));
    
    \ReadMemoryState[4]\ : SLE
      port map(D => ReadMemoryState_ns(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ReadMemoryState_Z(4));
    
    \mainProcess.pageaddr_5_i_m4[19]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(19), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(19), Y => N_4369);
    
    \mainProcess.InternalData2Memory_27_0_iv_3[13]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(13), B => 
        TimeStampValue(13), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_3(13));
    
    \StartAddrReg[26]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(26));
    
    \ControllUnitState_ns_i_0_1[11]\ : CFG4
      generic map(INIT => x"50DC")

      port map(A => N_4423, B => N_4339, C => dataReady_0, D => 
        ControllUnitState_Z(3), Y => 
        ControllUnitState_ns_i_0_1_Z(11));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[21]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(21), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0(21));
    
    InternalAddr2Memory_0_sqmuxa_2_i_a2_8 : CFG4
      generic map(INIT => x"4C00")

      port map(A => ControllUnitState_Z(4), B => 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_2_Z, C => N_4343_i, D
         => InternalAddr2Memory_0_sqmuxa_2_i_a2_6_Z, Y => 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_8_Z);
    
    \StampFSMR1[27]\ : SLE
      port map(D => pageaddr_5(27), CLK => sb_sb_0_FIC_0_CLK, EN
         => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(27));
    
    \mainProcess.PRDATA_8_0_iv_0[24]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(24), B => 
        PRDATA_8_0_iv_0_3(24), C => PRDATA_8_0_iv_0_6(24), Y => 
        PRDATA_8(24));
    
    \CommandReg[21]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(21));
    
    un1_memorycnt_1_s_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => memorycnt_Z(8), C => \GND\, D => 
        \GND\, FCI => un1_memorycnt_1_cry_7_Z, S => 
        un1_memorycnt_1_s_8_S, Y => un1_memorycnt_1_s_8_Y, FCO
         => un1_memorycnt_1_s_8_FCO);
    
    \mainProcess.PRDATA_8_0_iv_0_1[23]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize(15), B => CommandReg_Z(23), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(23));
    
    \StartAddrReg[31]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(31), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(31));
    
    \mainProcess.un1_readmemorycounter_0_o2\ : CFG4
      generic map(INIT => x"0010")

      port map(A => readmemorycounter_Z(3), B => 
        readmemorycounter_Z(2), C => readmemorycounter_Z(1), D
         => readmemorycounter_Z(0), Y => N_4272_i);
    
    un1_memorycnt_1_cry_1 : ARI1
      generic map(INIT => x"523DC")

      port map(A => memorycnt_Z(1), B => N_1260, C => 
        un23_0_0_Z(2), D => un23_0_a2_1_0_Z(2), FCI => \GND\, S
         => un1_memorycnt_1_cry_1_S, Y => un1_memorycnt_1_cry_1_Y, 
        FCO => un1_memorycnt_1_cry_1_Z);
    
    ControllUnitState_tr25_0_a2 : CFG4
      generic map(INIT => x"1000")

      port map(A => tempcounter_Z(2), B => tempcounter_Z(6), C
         => ControllUnitState_tr25_0_a2_5_Z, D => 
        ControllUnitState_tr25_0_a2_4_Z, Y => N_5700);
    
    \ConfigStatusReg[24]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(24));
    
    \ReadMemoryState_ns_i_0_a3[2]\ : CFG3
      generic map(INIT => x"31")

      port map(A => ReadMemoryState_Z(7), B => 
        ReadMemoryState_Z(6), C => N_68, Y => N_4286);
    
    \SPITransmitReg_RNO_0[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(0), Y => N_13_mux_1);
    
    \CommandReg[7]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(7));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[2]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(2), C => 
        Stamp1ShadowReg2_Z(2), D => 
        InternalData2Memory_27_0_iv_0_1(2), Y => 
        InternalData2Memory_27(2));
    
    \ReadMemoryState[8]\ : SLE
      port map(D => N_2471_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => ReadMemoryState_Z(8));
    
    \CurrentAddrReg[12]\ : SLE
      port map(D => un1_currentaddrreg_cry_12_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(12));
    
    Command_1_sqmuxa_0_a2_0_0 : CFG3
      generic map(INIT => x"04")

      port map(A => sb_sb_0_STAMP_PADDR(5), B => N_1025, C => 
        sb_sb_0_STAMP_PADDR(4), Y => Command_1_sqmuxa_0_a2_0_Z);
    
    \mainProcess.PRDATA_8_0_iv_0[30]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(30), B => 
        PRDATA_8_0_iv_0_3(30), C => PRDATA_8_0_iv_0_6(30), Y => 
        PRDATA_8(30));
    
    un1_readmemoryaddrcounter_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemoryaddrcounter_Z(27), C
         => \GND\, D => \GND\, FCI => 
        un1_readmemoryaddrcounter_cry_3_Z, S => 
        un1_readmemoryaddrcounter_cry_4_S, Y => 
        un1_readmemoryaddrcounter_cry_4_Y, FCO => 
        un1_readmemoryaddrcounter_cry_4_Z);
    
    \SPITransmitReg_RNO[28]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_3, B => InternalDataFromMem(28), C => 
        N_54, D => N_15_mux_2, Y => SPITransmitReg_13(28));
    
    \CommandReg[31]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(31), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(31));
    
    \CommandReg[14]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(14));
    
    \Stamp1ShadowReg2[14]\ : SLE
      port map(D => STAMP_0_data_frame(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(14));
    
    \mainProcess.PRDATA_8_0_iv_0[27]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(27), B => 
        PRDATA_8_0_iv_0_3(27), C => PRDATA_8_0_iv_0_6(27), Y => 
        PRDATA_8(27));
    
    \CommandReg[9]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(9));
    
    \Stamp1ShadowReg2[5]\ : SLE
      port map(D => STAMP_0_data_frame(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(5));
    
    \mainProcess.PRDATA_8_0_iv_0_3[8]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(8), B => 
        Stamp1ShadowReg2_Z(8), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(8));
    
    \SPITransmitReg_RNO_1[25]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(25), Y => N_15_mux_5);
    
    \Stamp1ShadowReg2[27]\ : SLE
      port map(D => STAMP_0_data_frame(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(27));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[10]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(10), C => 
        Stamp1ShadowReg2_Z(10), D => 
        InternalData2Memory_27_0_iv_0_1(10), Y => 
        InternalData2Memory_27(10));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[8]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(8), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(8));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[10]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(10), B => 
        TimeStampValue(10), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(10));
    
    \InternalData2Memory[2]\ : SLE
      port map(D => InternalData2Memory_27(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(2));
    
    \PRDATA[10]\ : SLE
      port map(D => PRDATA_8(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(10));
    
    \Command[1]\ : SLE
      port map(D => N_178_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        Command_1_sqmuxa_1_i_Z, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        Command_Z(1));
    
    WriteEnable_RNO : CFG4
      generic map(INIT => x"00BA")

      port map(A => ReadMemoryState_Z(4), B => 
        ReadMemoryState_Z(5), C => un1_ControllUnitState_9, D => 
        ReadMemoryState_ns(5), Y => N_4265_i);
    
    \readmemorycounter[3]\ : SLE
      port map(D => N_4262_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => readmemorycounter_Z(3));
    
    \un23_a3_1[1]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => ControllUnitState_Z(3), B => 
        ControllUnitSubState_Z(0), C => ControllUnitState_Z(5), D
         => ControllUnitState_Z(6), Y => N_1298);
    
    \mainProcess.PRDATA_8_0_iv_0_2[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(29), 
        D => CurrentAddrReg_Z(29), Y => PRDATA_8_0_iv_0_2(29));
    
    \readmemoryaddrcounter[26]\ : SLE
      port map(D => un1_readmemoryaddrcounter_cry_5_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemoryaddrcounter_Z(26));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[17]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(17), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(17));
    
    \CommandReg[11]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(11));
    
    \ReadMemoryState[7]\ : SLE
      port map(D => N_44, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryState_Z(7));
    
    \Stamp1ShadowReg2[23]\ : SLE
      port map(D => STAMP_0_data_frame(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(23));
    
    \SPITransmitReg_RNO_0[15]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(7), Y => N_4_16);
    
    \ConfigStatusReg[27]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(27));
    
    enableSPI_0_sqmuxa_2_0_a2_RNO : CFG3
      generic map(INIT => x"80")

      port map(A => counter_Z(1), B => InternalBusy, C => 
        counter_Z(0), Y => N_144);
    
    \ControllUnitSubState_RNIDU3L_0[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => ControllUnitSubState_Z(0), B => 
        ControllUnitSubState_Z(1), Y => N_4343_i);
    
    \SPIState[0]\ : SLE
      port map(D => N_154_mux_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \GND\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => SPIState_Z(0));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[3]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(3), C => 
        Stamp1ShadowReg2_Z(3), D => 
        InternalData2Memory_27_0_iv_0_1(3), Y => 
        InternalData2Memory_27(3));
    
    \mainProcess.InternalAddr2Memory_34_1[3]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => readmemorylimitedcnt_Z(3), B => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), C => N_138, Y
         => InternalAddr2Memory_34_1(3));
    
    \SPITransmitReg_RNO[10]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_21, B => InternalDataFromMem(10), C => 
        N_54, D => N_15_mux_20, Y => SPITransmitReg_13(10));
    
    \mainProcess.PRDATA_8_0_iv_0_0[8]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(8), D => SPIRecReg(8), Y => 
        PRDATA_8_0_iv_0_0(8));
    
    \mainProcess.pageaddr_5_i_m4[26]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(26), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(26), Y => pageaddr_5_i_m4(26));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[12]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(12), C => 
        Stamp1ShadowReg2_Z(12), D => 
        InternalData2Memory_27_0_iv_0_1(12), Y => 
        InternalData2Memory_27(12));
    
    \mainProcess.InternalAddr2Memory_34_1[5]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => readmemorylimitedcnt_Z(5), B => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), C => N_138, Y
         => InternalAddr2Memory_34_1(5));
    
    \MemoryPageSize[10]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(10));
    
    \mainProcess.PRDATA_8_0_iv_0_1[7]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ConfigStatusReg_Z(7), B => CommandReg_Z(7), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(7));
    
    \StampFSMPC[2]\ : SLE
      port map(D => StampFSMPC_6(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_1246_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => StampFSMPC_Z(2));
    
    \mainProcess.PRDATA_8_0_iv_0_1[11]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(3), B => CommandReg_Z(11), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(11));
    
    \ReadMemoryShadowReg[17]\ : SLE
      port map(D => InternalDataFromMem(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(17));
    
    \mainProcess.SPITransmitReg_13_0_iv_0[2]\ : CFG4
      generic map(INIT => x"A808")

      port map(A => N_4270, B => InternalDataFromMem(2), C => 
        SPIState_1_sqmuxa, D => sb_sb_0_STAMP_PWDATA(2), Y => 
        SPITransmitReg_13(2));
    
    \ReadMemoryShadowReg[21]\ : SLE
      port map(D => InternalDataFromMem(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(21));
    
    un1_currentaddrreg_cry_1 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize(1), B => pageaddr(1), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_0_Z, S
         => un1_currentaddrreg_cry_1_S, Y => 
        un1_currentaddrreg_cry_1_Y, FCO => 
        un1_currentaddrreg_cry_1_Z);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[15]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(15), B => 
        TimeStampValue(15), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(15));
    
    \SPITransmitReg_RNO_1[13]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(13), Y => N_15_mux_17);
    
    un1_currentaddrreg_cry_29 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(29), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_28_Z, S => 
        un1_currentaddrreg_cry_29_S, Y => 
        un1_currentaddrreg_cry_29_Y, FCO => 
        un1_currentaddrreg_cry_29_Z);
    
    \PRDATA[13]\ : SLE
      port map(D => PRDATA_8(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(13));
    
    \StampFSMPC_6_0_a2[2]\ : CFG2
      generic map(INIT => x"2")

      port map(A => un8_tempcounter_cry_2_S, B => 
        ControllUnitState_Z(11), Y => StampFSMPC_6(2));
    
    \CurrentAddrReg[29]\ : SLE
      port map(D => un1_currentaddrreg_cry_29_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(29));
    
    \ReadMemoryState_ns_i_o4_3[0]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => Command_Z(7), B => Command_Z(3), C => 
        Command_Z(2), D => Command_Z(1), Y => 
        ReadMemoryState_ns_i_o4_3_Z(0));
    
    \readmemorycounter_RNO[0]\ : CFG3
      generic map(INIT => x"2C")

      port map(A => N_1508_i, B => un1_enableSPI_1_sqmuxa_1_i, C
         => readmemorycounter_Z(0), Y => N_4260_i);
    
    \mainProcess.PRDATA_8_0_iv_0_2[0]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(0), 
        D => CurrentAddrReg_Z(0), Y => PRDATA_8_0_iv_0_2(0));
    
    \mainProcess.PRDATA_8_0_iv_0_0[16]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(16), D => SPIRecReg(16), Y => 
        PRDATA_8_0_iv_0_0(16));
    
    un1_SPIState_8_0_0 : CFG4
      generic map(INIT => x"FF2E")

      port map(A => SPIState_Z(3), B => N_62, C => N_4272_i, D
         => N_102, Y => un1_SPIState_8);
    
    \SPITransmitReg_RNO_1[29]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(29), Y => N_15_mux_1);
    
    \InternalAddr2Memory[2]\ : SLE
      port map(D => InternalAddr2Memory_34(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => InternalAddr2Memory_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => InternalAddr2Memory_Z(2));
    
    \ConfigStatusReg[7]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(7));
    
    \ConfigStatusReg[28]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(28));
    
    \Stamp1ShadowReg2[26]\ : SLE
      port map(D => STAMP_0_data_frame(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(26));
    
    \ConfigStatusReg_RNO[29]\ : CFG4
      generic map(INIT => x"0415")

      port map(A => SPIState_Z(1), B => SPIState_Z(3), C => 
        SPIState_ns(3), D => m98_xx_mm_1, Y => 
        ConfigStatusReg_40(29));
    
    \StartAddrReg[24]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(24));
    
    \ControllUnitState[7]\ : SLE
      port map(D => ControllUnitState_ns(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(7));
    
    \Command_RNO[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => sb_sb_0_STAMP_PWDATA(27), B => 
        SPIState_RNI27U44_Z(1), Y => N_174_i);
    
    \SPITransmitReg_RNO_1[22]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(22), Y => N_15_mux_8);
    
    \PRDATA[3]\ : SLE
      port map(D => PRDATA_8(3), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(3));
    
    \mainProcess.PRDATA_8_0_iv_0_6[3]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(3), C => 
        PRDATA_8_0_iv_0_1(3), D => PRDATA_8_0_iv_0_0(3), Y => 
        PRDATA_8_0_iv_0_6(3));
    
    \mainProcess.PRDATA_8_0_iv_0_1[24]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ConfigStatusReg_Z(24), B => CommandReg_Z(24), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(24));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[16]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(16), C => pageaddr(24), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(16));
    
    \InternalData2Memory[23]\ : SLE
      port map(D => InternalData2Memory_27(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(23));
    
    \ControllUnitSubState_ns_0_0_a2_0[0]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => N_2648, B => N_2631, C => N_1035, D => 
        enableSPI_1_sqmuxa_1_0_Z, Y => N_4614);
    
    \mainProcess.readmemorylimitedcnt_5[4]\ : CFG2
      generic map(INIT => x"2")

      port map(A => readmemorylimitedcnt_RNIBBFG2_S(4), B => 
        APB3ReadMemoryLimitedState_Z(1), Y => 
        readmemorylimitedcnt_5(4));
    
    \PRDATA[5]\ : SLE
      port map(D => PRDATA_8(5), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(5));
    
    un1_currentaddrreg_cry_3 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(3), B => pageaddr(3), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_2_Z, S
         => un1_currentaddrreg_cry_3_S, Y => 
        un1_currentaddrreg_cry_3_Y, FCO => 
        un1_currentaddrreg_cry_3_Z);
    
    \SPITransmitReg[18]\ : SLE
      port map(D => SPITransmitReg_13(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(18));
    
    \SPITransmitReg_RNO_0[19]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(11), Y => N_4_12);
    
    \mainProcess.PRDATA_8_0_iv_0_6[16]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(16), C => 
        PRDATA_8_0_iv_0_1(16), D => PRDATA_8_0_iv_0_0(16), Y => 
        PRDATA_8_0_iv_0_6(16));
    
    \SPITransmitReg_RNO_0[12]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(4), Y => N_4_19);
    
    \MemoryPageSize[6]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(6));
    
    \tempcounter[0]\ : SLE
      port map(D => tempcounter_7_iv_i(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_enabletimestampgen2_1_i, ALn
         => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, 
        LAT => \GND\, Q => tempcounter_Z(0));
    
    \SPIState_RNO_3[2]\ : CFG4
      generic map(INIT => x"0703")

      port map(A => Command_Z(0), B => SPIState_Z(4), C => 
        SPIState_ns(3), D => N_21_0, Y => N_150_mux);
    
    un1_enabletimestampgen2_5_3 : CFG4
      generic map(INIT => x"EEFE")

      port map(A => ControllUnitState_Z(0), B => 
        ControllUnitState_Z(1), C => ControllUnitState_Z(3), D
         => ControllUnitSubState_Z(0), Y => 
        un1_enabletimestampgen2_5_3_Z);
    
    \StartAddrReg[10]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(10));
    
    \mainProcess.PRDATA_8_0_iv_0_3[17]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(17), B => 
        Stamp1ShadowReg2_Z(17), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(17));
    
    \StampFSMPC[7]\ : SLE
      port map(D => StampFSMPC_6(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_1246_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => StampFSMPC_Z(7));
    
    \InternalData2Memory[25]\ : SLE
      port map(D => InternalData2Memory_27(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(25));
    
    \mainProcess.InternalData2Memory_27_0_iv[11]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_3(11), C => 
        Stamp1ShadowReg2_Z(11), D => 
        InternalData2Memory_27_0_iv_1(11), Y => 
        InternalData2Memory_27(11));
    
    \mainProcess.pageaddr_5_i_m4[25]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(25), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(25), Y => pageaddr_5_i_m4(25));
    
    \StampFSMPC_6[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => un8_tempcounter_cry_1_S, B => 
        ControllUnitState_Z(11), Y => StampFSMPC_6_Z(1));
    
    \ReadMemoryShadowReg[20]\ : SLE
      port map(D => InternalDataFromMem(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(20));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[6]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(6), C => 
        Stamp1ShadowReg2_Z(6), D => 
        InternalData2Memory_27_0_iv_0_1(6), Y => 
        InternalData2Memory_27(6));
    
    \APB3ReadMemoryLimitedState_RNI12J4[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => APB3ReadMemoryLimitedState_Z(5), 
        C => ConfigStatusReg_Z(4), D => \GND\, FCI => \VCC\, S
         => APB3ReadMemoryLimitedState_RNI12J4_S(5), Y => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), FCO => 
        un1_readmemorylimitedcnt_cry_0_cy);
    
    \SPITransmitReg_RNO[27]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_4, B => InternalDataFromMem(27), C => 
        N_54, D => N_15_mux_3, Y => SPITransmitReg_13(27));
    
    PREADY_1_i_a2_0_a4 : CFG2
      generic map(INIT => x"E")

      port map(A => APBState_Z(1), B => APBState_Z(0), Y => 
        N_1539_i);
    
    \mainProcess.PRDATA_8_0_iv_0_3[6]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(6), B => 
        Stamp1ShadowReg2_Z(6), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(6));
    
    \InternalAddr2Memory[4]\ : SLE
      port map(D => InternalAddr2Memory_34(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => InternalAddr2Memory_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => InternalAddr2Memory_Z(4));
    
    \Stamp1ShadowReg1[21]\ : SLE
      port map(D => STAMP_0_data_frame(53), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(21));
    
    \readmemoryaddrcounter[25]\ : SLE
      port map(D => un1_readmemoryaddrcounter_cry_6_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemoryaddrcounter_Z(25));
    
    \StampFSMPC[0]\ : SLE
      port map(D => N_746_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_1246_i, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => StampFSMPC_Z(0));
    
    \SPIState_RNO[0]\ : CFG4
      generic map(INIT => x"FF20")

      port map(A => N_154_mux_i_1_0, B => SPIState_1_sqmuxa, C
         => SPIState_Z(0), D => SPIState_Z(1), Y => N_154_mux_i);
    
    \MemoryPageSize[2]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(2));
    
    \mainProcess.SPIaddr_15_iv_0_m2_RNO[0]\ : CFG4
      generic map(INIT => x"C0E2")

      port map(A => ControllUnitState_Z(1), B => N_23_0, C => 
        Command_Z(4), D => SPIaddr_Z(0), Y => N_155_mux_i);
    
    \mainProcess.InternalAddr2Memory_34_1[6]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => readmemorylimitedcnt_Z(6), B => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), C => N_138, Y
         => InternalAddr2Memory_34_1(6));
    
    \mainProcess.PRDATA_8_0_iv_0_6[25]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(25), C => 
        PRDATA_8_0_iv_0_1(25), D => PRDATA_8_0_iv_0_0(25), Y => 
        PRDATA_8_0_iv_0_6(25));
    
    \Stamp1ShadowReg1[18]\ : SLE
      port map(D => STAMP_0_data_frame(50), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(18));
    
    un1_currentaddrreg_cry_27 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(27), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_26_Z, S => 
        un1_currentaddrreg_cry_27_S, Y => 
        un1_currentaddrreg_cry_27_Y, FCO => 
        un1_currentaddrreg_cry_27_Z);
    
    \SPITransmitReg[25]\ : SLE
      port map(D => SPITransmitReg_13(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(25));
    
    \mainProcess.readmemorylimitedcnt_5[6]\ : CFG2
      generic map(INIT => x"2")

      port map(A => readmemorylimitedcnt_RNIMSQE3_S(6), B => 
        APB3ReadMemoryLimitedState_Z(1), Y => 
        readmemorylimitedcnt_5(6));
    
    \ConfigStatusReg_RNO_3[4]\ : CFG3
      generic map(INIT => x"04")

      port map(A => APB3ReadMemoryLimitedState_Z(1), B => 
        m84_m7_0, C => sb_sb_0_STAMP_PADDR(11), Y => m84_m7_1);
    
    \APBState_RNIA9JC[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => ReadMemoryState_Z(3), B => APBState_Z(1), Y
         => m84_m7_0);
    
    \InternalData2Memory[8]\ : SLE
      port map(D => InternalData2Memory_27(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(8));
    
    \CurrentAddrReg[3]\ : SLE
      port map(D => un1_currentaddrreg_cry_3_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(3));
    
    \ReadMemoryShadowReg[24]\ : SLE
      port map(D => InternalDataFromMem(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(24));
    
    \ConfigStatusReg_RNO[4]\ : CFG3
      generic map(INIT => x"87")

      port map(A => m84_N_13_mux, B => r_N_6_mux, C => d_N_5_mux, 
        Y => N_85_i);
    
    \un23_0_a2_1_0[2]\ : CFG4
      generic map(INIT => x"1110")

      port map(A => ControllUnitState_Z(8), B => 
        ControllUnitState_Z(6), C => ControllUnitSubState_Z(1), D
         => ControllUnitSubState_Z(0), Y => un23_0_a2_1_0_Z(2));
    
    \ReadMemoryState_RNO[6]\ : CFG4
      generic map(INIT => x"0A08")

      port map(A => N_4274, B => ReadMemoryState_Z(7), C => 
        N_4286, D => N_2496, Y => N_2475_i);
    
    \memorycnt[2]\ : SLE
      port map(D => memorycnt_6(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => memorycnt_Z(2));
    
    \mainProcess.SPIaddr_15_iv_0_RNO[0]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => SPIaddr_0_sqmuxa_3, B => isfirstrun_Z(0), C
         => ControllUnitState_RNI2VHT_Z(14), D => N_23_0, Y => 
        SPIaddr_3_sqmuxa_1);
    
    \CurrentAddrReg[5]\ : SLE
      port map(D => un1_currentaddrreg_cry_5_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(5));
    
    un1_memorycnt_1_cry_2 : ARI1
      generic map(INIT => x"513EC")

      port map(A => memorycnt_Z(2), B => N_1262, C => un23_1_Z(1), 
        D => un23_a3_0(1), FCI => un1_memorycnt_1_cry_1_Z, S => 
        un1_memorycnt_1_cry_2_S, Y => un1_memorycnt_1_cry_2_Y, 
        FCO => un1_memorycnt_1_cry_2_Z);
    
    \SPITransmitReg_RNO[22]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_9, B => InternalDataFromMem(22), C => 
        N_54, D => N_15_mux_8, Y => SPITransmitReg_13(22));
    
    \ControllUnitState_RNI2VHT_0[14]\ : CFG1
      generic map(INIT => "01")

      port map(A => ControllUnitState_RNI2VHT_Z(14), Y => 
        N_1541_i);
    
    \CommandReg[5]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(5));
    
    un1_memorycnt_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => memorycnt_Z(6), C => \GND\, D => 
        \GND\, FCI => un1_memorycnt_1_cry_5_Z, S => 
        un1_memorycnt_1_cry_6_S, Y => un1_memorycnt_1_cry_6_Y, 
        FCO => un1_memorycnt_1_cry_6_Z);
    
    \SPIState_RNO[3]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => Command_Z(0), B => SPIState_Z(4), C => 
        N_2496_i, D => N_21_0, Y => N_70);
    
    \ReadMemoryShadowReg[19]\ : SLE
      port map(D => InternalDataFromMem(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(19));
    
    \mainProcess.PRDATA_8_0_iv_0_0[18]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(18), D => SPIRecReg(18), Y => 
        PRDATA_8_0_iv_0_0(18));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[22]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(22), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(22));
    
    \SPIState_RNO_0[2]\ : CFG4
      generic map(INIT => x"4C0C")

      port map(A => SPIState_Z(4), B => SPIState_Z(2), C => 
        m41_0_2_1, D => SPIState_1_sqmuxa, Y => m41_0_1);
    
    \mainProcess.pageaddr_5_i_m4[20]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(20), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(20), Y => pageaddr_5_i_m4(20));
    
    \APB3ReadMemoryLimitedState[4]\ : SLE
      port map(D => APB3ReadMemoryLimitedState_RNI12J4_Y(5), CLK
         => sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => APB3ReadMemoryLimitedState_Z(4));
    
    enableSPI_1_sqmuxa_1_0 : CFG2
      generic map(INIT => x"8")

      port map(A => ControllUnitState_Z(2), B => 
        ControllUnitSubState_Z(1), Y => enableSPI_1_sqmuxa_1_0_Z);
    
    \Command_RNI6AH02_0[1]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => Command_Z(1), B => m17_e_1, C => Command_Z(3), 
        D => Command_Z(2), Y => N_19_0);
    
    \mainProcess.PRDATA_8_0_iv_0_0[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(29), D => SPIRecReg(29), Y => 
        PRDATA_8_0_iv_0_0(29));
    
    \mainProcess.pageaddr_5_i_m4[24]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(24), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(24), Y => pageaddr_5_i_m4(24));
    
    \mainProcess.InternalAddr2Memory_34[2]\ : CFG4
      generic map(INIT => x"FDDD")

      port map(A => InternalAddr2Memory_34_1(2), B => 
        InternalAddr2Memory_34_18, C => 
        readmemoryaddrcounter_Z(29), D => ReadMemoryState_Z(4), Y
         => InternalAddr2Memory_34(2));
    
    \ConfigStatusReg[9]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize(1));
    
    \SPITransmitReg_RNO[16]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_15, B => InternalDataFromMem(16), C => 
        N_54, D => N_15_mux_14, Y => SPITransmitReg_13(16));
    
    \PRDATA[15]\ : SLE
      port map(D => PRDATA_8(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(15));
    
    \mainProcess.InternalAddr2Memory_34_22\ : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory_34_sm0, B => 
        InternalAddr2Memory_34_m0(6), C => N_143_mux, Y => 
        InternalAddr2Memory_34_22);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[14]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(14), B => 
        TimeStampValue(14), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(14));
    
    un1_currentaddrreg_cry_11 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(11), B => pageaddr(11), C
         => \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_10_Z, 
        S => un1_currentaddrreg_cry_11_S, Y => 
        un1_currentaddrreg_cry_11_Y, FCO => 
        un1_currentaddrreg_cry_11_Z);
    
    \PRDATA[6]\ : SLE
      port map(D => PRDATA_8(6), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(6));
    
    \mainProcess.PRDATA_8_0_iv_0_6[31]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(31), C => 
        PRDATA_8_0_iv_0_1(31), D => PRDATA_8_0_iv_0_0(31), Y => 
        PRDATA_8_0_iv_0_6(31));
    
    \SPIState_RNI54C35[4]\ : CFG4
      generic map(INIT => x"F838")

      port map(A => N_19_0, B => SPIState_Z(4), C => m106_1_1, D
         => N_21_0, Y => N_23_0);
    
    \mainProcess.PRDATA_8_0_iv_0_2[6]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(6), 
        D => CurrentAddrReg_Z(6), Y => PRDATA_8_0_iv_0_2(6));
    
    \MemoryPageSize[13]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(13));
    
    \mainProcess.PRDATA_8_0_iv_0_6[18]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(18), C => 
        PRDATA_8_0_iv_0_1(18), D => PRDATA_8_0_iv_0_0(18), Y => 
        PRDATA_8_0_iv_0_6(18));
    
    \counter[0]\ : SLE
      port map(D => N_140_mux_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => counter_Z(0));
    
    \CommandReg[26]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(26));
    
    \Stamp1ShadowReg1[7]\ : SLE
      port map(D => STAMP_0_data_frame(39), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(7));
    
    \ConfigStatusReg[4]\ : SLE
      port map(D => N_85_i, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ConfigStatusReg_Z(4));
    
    un1_readmemoryaddrcounter_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemoryaddrcounter_Z(30), C
         => \GND\, D => \GND\, FCI => 
        un1_readmemoryaddrcounter_cry_0_Z, S => 
        un1_readmemoryaddrcounter_cry_1_S, Y => 
        un1_readmemoryaddrcounter_cry_1_Y, FCO => 
        un1_readmemoryaddrcounter_cry_1_Z);
    
    \StampFSMR1[7]\ : SLE
      port map(D => pageaddr_5_i_m4(7), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(7));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[20]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(20), B => 
        TimeStampValue(20), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(20));
    
    InternalAddr2Memory_0_sqmuxa_2_i_a2_6 : CFG4
      generic map(INIT => x"3050")

      port map(A => ControllUnitState_Z(2), B => 
        ControllUnitState_Z(6), C => N_1128, D => N_4343_i, Y => 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_6_Z);
    
    \ControllUnitSubState_ns_0_0_o4[0]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => ConfigStatusReg_Z(2), B => 
        ControllUnitState_Z(0), C => N_2631, D => N_1035, Y => 
        N_4346);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[3]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(3), C => pageaddr(11), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(3));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[8]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(8), C => 
        Stamp1ShadowReg2_Z(8), D => 
        InternalData2Memory_27_0_iv_0_1(8), Y => 
        InternalData2Memory_27(8));
    
    InternalAddr2Memory_11_sqmuxa_i_o3 : CFG2
      generic map(INIT => x"7")

      port map(A => GPIO_6_M2F_c, B => ControllUnitSubState_Z(0), 
        Y => N_1255_i);
    
    \mainProcess.PRDATA_8_0_iv_0_2[17]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(17), 
        D => CurrentAddrReg_Z(17), Y => PRDATA_8_0_iv_0_2(17));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_a2_1[23]\ : CFG3
      generic map(INIT => x"02")

      port map(A => TimeStampValue(23), B => ReadMemoryState_Z(4), 
        C => N_1232_i, Y => N_4527);
    
    \counter_RNIG30C1[0]\ : CFG3
      generic map(INIT => x"20")

      port map(A => counter_Z(1), B => InternalBusy, C => 
        counter_Z(0), Y => counter9);
    
    \ControllUnitState[1]\ : SLE
      port map(D => ControllUnitState_ns(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(1));
    
    \SPITransmitReg[27]\ : SLE
      port map(D => SPITransmitReg_13(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(27));
    
    \mainProcess.PRDATA_8_0_iv_0[13]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(13), B => 
        PRDATA_8_0_iv_0_3(13), C => PRDATA_8_0_iv_0_6(13), Y => 
        PRDATA_8(13));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[20]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(20), C => 
        Stamp1ShadowReg2_Z(20), D => 
        InternalData2Memory_27_0_iv_0_1(20), Y => 
        InternalData2Memory_27(20));
    
    \ControllUnitSubState[1]\ : SLE
      port map(D => N_2629_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        GPIO_6_M2F_c, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ControllUnitSubState_Z(1));
    
    \mainProcess.PRDATA_8_0_iv_0[22]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(22), B => 
        PRDATA_8_0_iv_0_3(22), C => PRDATA_8_0_iv_0_6(22), Y => 
        PRDATA_8(22));
    
    \mainProcess.InternalData2Memory_27_0_iv_3[21]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(21), B => 
        TimeStampValue(21), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_3(21));
    
    \ControllUnitState_ns_0_a5_0_a2[13]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_4353, B => ControllUnitState_Z(2), Y => 
        ControllUnitState_ns(13));
    
    \tempcounter_RNO[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_1261_i, B => un8_tempcounter_cry_1_S, Y => 
        tempcounter_7(1));
    
    \StartAddrReg[9]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(9));
    
    \mainProcess.InternalAddr2Memory_34_m4_0[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => ReadMemoryState_Z(4), B => 
        readmemoryaddrcounter_Z(30), Y => 
        InternalAddr2Memory_34_m4(1));
    
    InternalAddr2Memory_0_sqmuxa_2_i_a2_2 : CFG3
      generic map(INIT => x"D0")

      port map(A => ControllUnitState_Z(3), B => 
        ControllUnitSubState_Z(0), C => 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_1_Z, Y => 
        InternalAddr2Memory_0_sqmuxa_2_i_a2_2_Z);
    
    SPIaddr_2_sqmuxa_1_i_0 : CFG4
      generic map(INIT => x"AEFF")

      port map(A => N_23_0, B => GPIO_6_M2F_c, C => N_4424, D => 
        SPIaddr_0_sqmuxa_3, Y => N_127);
    
    \ReadMemoryState_RNIKQ802[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => SPIState_ns(3), B => ReadMemoryState_Z(3), Y
         => SPIaddr_0_sqmuxa_3);
    
    \mainProcess.PRDATA_8_0_iv_0_1[1]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ConfigStatusReg_Z(1), B => CommandReg_Z(1), C
         => N_1025, D => N_4335, Y => PRDATA_8_0_iv_0_1(1));
    
    \mainProcess.PRDATA_8_0_iv_0_2[26]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(26), 
        D => CurrentAddrReg_Z(26), Y => PRDATA_8_0_iv_0_2(26));
    
    \mainProcess.un1_paddr_3\ : CFG3
      generic map(INIT => x"04")

      port map(A => sb_sb_0_STAMP_PADDR(2), B => 
        sb_sb_0_STAMP_PADDR(6), C => sb_sb_0_STAMP_PADDR(3), Y
         => un1_paddr_3);
    
    \readmemorycounter[2]\ : SLE
      port map(D => N_4261_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => readmemorycounter_Z(2));
    
    \Stamp1ShadowReg1[24]\ : SLE
      port map(D => STAMP_0_data_frame(56), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(24));
    
    \APB3ReadMemoryLimitedState_RNO_0[0]\ : CFG4
      generic map(INIT => x"51FB")

      port map(A => APB3ReadMemoryLimitedState_Z(0), B => 
        ConfigStatusReg_Z(4), C => 
        APB3ReadMemoryLimitedState_Z(1), D => PRDATA_17_sqmuxa_Z, 
        Y => N_50_0);
    
    Command_1_sqmuxa_0_a2 : CFG4
      generic map(INIT => x"0400")

      port map(A => sb_sb_0_STAMP_PADDR(11), B => 
        Command_1_sqmuxa_0_a2_1_0_Z, C => un1_APBState_1_2_0_Z, D
         => Command_1_sqmuxa_0_a2_0_Z, Y => Command_1_sqmuxa);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[17]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(17), C => pageaddr(25), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(17));
    
    \Stamp1ShadowReg2[21]\ : SLE
      port map(D => STAMP_0_data_frame(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(21));
    
    \CommandReg[16]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(16));
    
    \ReadMemoryShadowReg[22]\ : SLE
      port map(D => InternalDataFromMem(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(22));
    
    \MemoryPageSize[9]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \GND\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(9));
    
    \StartAddrReg[22]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(22));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[22]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(22), C => 
        Stamp1ShadowReg2_Z(22), D => 
        InternalData2Memory_27_0_iv_0_1(22), Y => 
        InternalData2Memory_27(22));
    
    \memorycnt[8]\ : SLE
      port map(D => memorycnt_6(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => memorycnt_Z(8));
    
    \mainProcess.InternalAddr2Memory_34_m5[1]\ : CFG4
      generic map(INIT => x"88F0")

      port map(A => readmemorylimitedcnt_Z(1), B => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), C => 
        InternalAddr2Memory_34_m4(1), D => N_138, Y => 
        InternalAddr2Memory_34_m5(1));
    
    \StartAddrReg[0]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(0));
    
    \ReadMemoryState[6]\ : SLE
      port map(D => N_2475_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => ReadMemoryState_Z(6));
    
    SPIState_m2_e_1_0 : CFG3
      generic map(INIT => x"7F")

      port map(A => sb_sb_0_STAMP_PADDR(4), B => 
        sb_sb_0_STAMP_PADDR(3), C => sb_sb_0_STAMP_PADDR(2), Y
         => SPIState_m2_e_1_0_Z);
    
    \SPITransmitReg_RNO_1[23]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(23), Y => N_15_mux_7);
    
    \SPITransmitReg[21]\ : SLE
      port map(D => SPITransmitReg_13(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(21));
    
    \Stamp1ShadowReg2[1]\ : SLE
      port map(D => STAMP_0_data_frame(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(1));
    
    \un23_i_a2[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => ControllUnitState_Z(4), B => 
        ControllUnitSubState_Z(0), C => ControllUnitState_Z(5), D
         => ControllUnitState_Z(6), Y => N_761);
    
    \StampFSMPC_6_0_a2[8]\ : CFG2
      generic map(INIT => x"2")

      port map(A => un8_tempcounter_s_8_S, B => 
        ControllUnitState_Z(11), Y => StampFSMPC_6(8));
    
    \mainProcess.PRDATA_8_0_iv_0_0[11]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(11), D => SPIRecReg(11), Y => 
        PRDATA_8_0_iv_0_0(11));
    
    \mainProcess.PRDATA_8_0_iv_0[11]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(11), B => 
        PRDATA_8_0_iv_0_3(11), C => PRDATA_8_0_iv_0_6(11), Y => 
        PRDATA_8(11));
    
    \CurrentAddrReg[4]\ : SLE
      port map(D => un1_currentaddrreg_cry_4_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(4));
    
    \mainProcess.InternalAddr2Memory_34_m2_1_1[1]\ : CFG3
      generic map(INIT => x"51")

      port map(A => ControllUnitState_Z(11), B => StampFSMPC_Z(1), 
        C => ControllUnitState_Z(10), Y => 
        InternalAddr2Memory_34_m2_1_1(1));
    
    un1_enabletimestampgen2_7_0_a3 : CFG3
      generic map(INIT => x"10")

      port map(A => ControllUnitState_Z(3), B => 
        ControllUnitState_Z(11), C => N_1254, Y => N_1302);
    
    \Stamp1ShadowReg1[9]\ : SLE
      port map(D => STAMP_0_data_frame(41), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(9));
    
    \mainProcess.PRDATA_8_0_iv_0_6[20]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(20), C => 
        PRDATA_8_0_iv_0_1(20), D => PRDATA_8_0_iv_0_0(20), Y => 
        PRDATA_8_0_iv_0_6(20));
    
    \InternalData2Memory[0]\ : SLE
      port map(D => InternalData2Memory_27(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(0));
    
    \ControllUnitState[9]\ : SLE
      port map(D => ControllUnitState_ns(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(9));
    
    \Stamp1ShadowReg2[18]\ : SLE
      port map(D => STAMP_0_data_frame(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(18));
    
    \mainProcess.ConfigStatusReg_26_0_a2_1[30]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => ControllUnitState_Z(3), B => dataReady_0, C
         => ConfigStatusReg_24_sn_N_11_mux, D => GPIO_6_M2F_c, Y
         => ConfigStatusReg_26_0_a2_1(30));
    
    \mainProcess.InternalAddr2Memory_34[6]\ : CFG4
      generic map(INIT => x"FDDD")

      port map(A => InternalAddr2Memory_34_1(6), B => 
        InternalAddr2Memory_34_22, C => 
        readmemoryaddrcounter_Z(25), D => ReadMemoryState_Z(4), Y
         => InternalAddr2Memory_34(6));
    
    \mainProcess.PRDATA_8_0_iv_0_6[5]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(5), C => 
        PRDATA_8_0_iv_0_1(5), D => PRDATA_8_0_iv_0_0(5), Y => 
        PRDATA_8_0_iv_0_6(5));
    
    \SPITransmitReg_RNO[11]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_20, B => InternalDataFromMem(11), C => 
        N_54, D => N_15_mux_19, Y => SPITransmitReg_13(11));
    
    \PRDATA[12]\ : SLE
      port map(D => PRDATA_8(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(12));
    
    \StartAddrReg[23]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(23));
    
    \ReadMemoryState_ns_i_0_0[3]\ : CFG4
      generic map(INIT => x"A0B3")

      port map(A => ReadMemoryState_ns_i_0_a3_2_8_Z(3), B => N_68, 
        C => ReadMemoryState_ns_i_0_a3_2_7_Z(3), D => 
        ReadMemoryState_Z(4), Y => ReadMemoryState_ns_i_0_0_Z(3));
    
    InternalData2Memory_5_sqmuxa : CFG3
      generic map(INIT => x"04")

      port map(A => N_1257_i, B => ControllUnitState_Z(9), C => 
        ReadMemoryState_Z(4), Y => InternalData2Memory_5_sqmuxa_Z);
    
    \mainProcess.readmemorycounter_6_iv_RNO_0[1]\ : CFG3
      generic map(INIT => x"80")

      port map(A => InternalBusy, B => N_62, C => N_4272_i, Y => 
        N_4254_i);
    
    un8_tempcounter_s_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => StampFSMPC_Z(8), C => \GND\, D
         => \GND\, FCI => un8_tempcounter_cry_7_Z, S => 
        un8_tempcounter_s_8_S, Y => un8_tempcounter_s_8_Y, FCO
         => un8_tempcounter_s_8_FCO);
    
    \ControllUnitSubState_ns_0_o2[0]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => ControllUnitState_Z(14), B => 
        ControllUnitState_Z(11), C => ControllUnitState_Z(13), Y
         => N_2631);
    
    \InternalData2Memory[28]\ : SLE
      port map(D => InternalData2Memory_27(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(28));
    
    \mainProcess.PRDATA_8_0_iv_0[15]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(15), B => 
        PRDATA_8_0_iv_0_3(15), C => PRDATA_8_0_iv_0_6(15), Y => 
        PRDATA_8(15));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[18]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(18), B => 
        TimeStampValue(18), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(18));
    
    \CurrentAddrReg[18]\ : SLE
      port map(D => un1_currentaddrreg_cry_18_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(18));
    
    \SPITransmitReg_RNO_0[13]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(5), Y => N_4_18);
    
    \SPIState_RNO[2]\ : CFG4
      generic map(INIT => x"0023")

      port map(A => SPIState_Z(3), B => SPIState_Z(1), C => 
        m41_0_1, D => SPIState_RNO_1_Z(2), Y => N_42_0);
    
    \PRDATA[19]\ : SLE
      port map(D => PRDATA_8(19), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(19));
    
    \mainProcess.pageaddr_5_i_m4[30]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(30), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(30), Y => pageaddr_5_i_m4(30));
    
    \ReadMemoryShadowReg[28]\ : SLE
      port map(D => InternalDataFromMem(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(28));
    
    un8_tempcounter_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => StampFSMPC_Z(3), C => \GND\, D
         => \GND\, FCI => un8_tempcounter_cry_2_Z, S => 
        un8_tempcounter_cry_3_S, Y => un8_tempcounter_cry_3_Y, 
        FCO => un8_tempcounter_cry_3_Z);
    
    \CurrentAddrReg[13]\ : SLE
      port map(D => un1_currentaddrreg_cry_13_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(13));
    
    \ControllUnitSubState_ns_0_0[0]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => N_1185, B => 
        ControllUnitSubState_ns_0_0_a2_1_Z(0), C => N_4346, D => 
        N_4614, Y => ControllUnitSubState_ns(0));
    
    \mainProcess.PRDATA_8_0_iv_0_6[11]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(11), C => 
        PRDATA_8_0_iv_0_1(11), D => PRDATA_8_0_iv_0_0(11), Y => 
        PRDATA_8_0_iv_0_6(11));
    
    un1_currentaddrreg_cry_19 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(19), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_18_Z, S => 
        un1_currentaddrreg_cry_19_S, Y => 
        un1_currentaddrreg_cry_19_Y, FCO => 
        un1_currentaddrreg_cry_19_Z);
    
    \ReadMemoryState_ns_i_0_o2[2]\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => readmemorycounter_Z(3), B => 
        readmemorycounter_Z(2), C => readmemorycounter_Z(1), D
         => readmemorycounter_Z(0), Y => N_4274);
    
    \mainProcess.PRDATA_8_0_iv_0_6[22]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(22), C => 
        PRDATA_8_0_iv_0_1(22), D => PRDATA_8_0_iv_0_0(22), Y => 
        PRDATA_8_0_iv_0_6(22));
    
    \ConfigStatusReg_RNO_0[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => sb_sb_0_STAMP_PADDR(7), B => 
        sb_sb_0_STAMP_PADDR(10), C => ConfigStatusReg_RNO_2_Z(4), 
        D => m84_m7_1, Y => m84_N_13_mux);
    
    \SPITransmitReg_RNO_0[28]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(20), Y => N_4_3);
    
    \ControllUnitSubState_ns_i_a7_4_4[1]\ : CFG3
      generic map(INIT => x"10")

      port map(A => memorycnt_Z(6), B => memorycnt_Z(5), C => 
        N_2624_1, Y => ControllUnitSubState_ns_i_a7_4_4_Z(1));
    
    \ConfigStatusReg_RNO_2[4]\ : CFG3
      generic map(INIT => x"A6")

      port map(A => N_81, B => sb_sb_0_STAMP_PWDATA(4), C => 
        N_2496_i, Y => ConfigStatusReg_RNO_2_Z(4));
    
    \ReadMemoryShadowReg[0]\ : SLE
      port map(D => InternalDataFromMem(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(0));
    
    \mainProcess.PRDATA_8_0_iv_0_6[23]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(23), C => 
        PRDATA_8_0_iv_0_1(23), D => PRDATA_8_0_iv_0_0(23), Y => 
        PRDATA_8_0_iv_0_6(23));
    
    \mainProcess.memorycnt_6_s_7\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => N_1541_i, C => memorycnt_Z(8), D
         => \GND\, FCI => memorycnt_6_cry_6, S => memorycnt_6(8), 
        Y => memorycnt_6_s_7_Y, FCO => memorycnt_6_s_7_FCO);
    
    ControllUnitSubState_2_sqmuxa_i_o3 : CFG3
      generic map(INIT => x"DF")

      port map(A => ControllUnitState_Z(2), B => N_5700, C => 
        ControllUnitSubState_Z(0), Y => N_1261_i);
    
    \SPITransmitReg[14]\ : SLE
      port map(D => SPITransmitReg_13(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(14));
    
    \SPITransmitReg[12]\ : SLE
      port map(D => SPITransmitReg_13(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(12));
    
    \mainProcess.PRDATA_8_0_iv_0_2[2]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(2), 
        D => CurrentAddrReg_Z(2), Y => PRDATA_8_0_iv_0_2(2));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[19]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(19), B => 
        TimeStampValue(19), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(19));
    
    \ConfigStatusReg_RNO[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => sb_sb_0_STAMP_PWDATA(31), B => N_4347, C => 
        N_4340, Y => N_249_i);
    
    \ReadMemoryShadowReg[9]\ : SLE
      port map(D => InternalDataFromMem(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(9));
    
    \Command[6]\ : SLE
      port map(D => N_168_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        Command_1_sqmuxa_1_i_Z, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        Command_Z(6));
    
    \StartAddrReg[16]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(16));
    
    \tempcounter[1]\ : SLE
      port map(D => tempcounter_7(1), CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_enabletimestampgen2_1_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => tempcounter_Z(1));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[5]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(5), B => TimeStampValue(5), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(5));
    
    \mainProcess.readmemorycounter_6_iv_RNO[1]\ : CFG4
      generic map(INIT => x"D31F")

      port map(A => N_1508_i, B => un1_enableSPI_1_sqmuxa_1_i, C
         => readmemorycounter_Z(1), D => readmemorycounter_Z(0), 
        Y => N_4259);
    
    \mainProcess.PRDATA_8_0_iv_0_3[27]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(27), B => 
        Stamp1ShadowReg2_Z(27), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(27));
    
    \mainProcess.PRDATA_8_0_iv_0_2[28]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(28), 
        D => CurrentAddrReg_Z(28), Y => PRDATA_8_0_iv_0_2(28));
    
    \mainProcess.memorycnt_6_cry_3\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => N_1541_i, C => memorycnt_Z(4), D
         => \GND\, FCI => memorycnt_6_cry_2, S => memorycnt_6(4), 
        Y => memorycnt_6_cry_3_Y, FCO => memorycnt_6_cry_3);
    
    \SPIState_RNO_2[2]\ : CFG4
      generic map(INIT => x"0F01")

      port map(A => SPIState_Z(4), B => m33_e_0, C => counter9, D
         => SPIState_RNO_5_Z(2), Y => m41_0_2_1);
    
    \StartAddrReg[30]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(30));
    
    \Command_RNO[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => sb_sb_0_STAMP_PWDATA(24), B => 
        SPIState_RNI27U44_Z(1), Y => N_180_i);
    
    \ControllUnitState_ns_i_a2_3[11]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => memorycnt_Z(6), B => memorycnt_Z(5), C => 
        memorycnt_Z(3), D => N_2624_2, Y => 
        ControllUnitState_ns_i_a2_3_Z(11));
    
    \mainProcess.PRDATA_8_0_iv_0_a2_9[12]\ : CFG3
      generic map(INIT => x"80")

      port map(A => sb_sb_0_STAMP_PADDR(2), B => 
        sb_sb_0_STAMP_PADDR(6), C => sb_sb_0_STAMP_PADDR(3), Y
         => N_1031);
    
    \mainProcess.PRDATA_8_0_iv_0[6]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(6), B => 
        PRDATA_8_0_iv_0_3(6), C => PRDATA_8_0_iv_0_6(6), Y => 
        PRDATA_8(6));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[9]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(9), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(9));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[10]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(10), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(10));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[16]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(16), C => 
        Stamp1ShadowReg2_Z(16), D => 
        InternalData2Memory_27_0_iv_0_1(16), Y => 
        InternalData2Memory_27(16));
    
    un1_APBState_1_1_0_a2_2 : CFG3
      generic map(INIT => x"01")

      port map(A => sb_sb_0_STAMP_PADDR(3), B => 
        sb_sb_0_STAMP_PADDR(5), C => sb_sb_0_STAMP_PADDR(4), Y
         => N_1028);
    
    \PRDATA[21]\ : SLE
      port map(D => PRDATA_8(21), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(21));
    
    \StampFSMR1[16]\ : SLE
      port map(D => pageaddr_5_i_m4(16), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(16));
    
    \Command_RNO[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => sb_sb_0_STAMP_PWDATA(29), B => 
        SPIState_RNI27U44_Z(1), Y => N_170_i);
    
    \SPITransmitReg[1]\ : SLE
      port map(D => SPITransmitReg_13(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(1));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[17]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(17), C => 
        Stamp1ShadowReg2_Z(17), D => 
        InternalData2Memory_27_0_iv_0_1(17), Y => 
        InternalData2Memory_27(17));
    
    \InternalData2Memory[11]\ : SLE
      port map(D => InternalData2Memory_27(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(11));
    
    \readmemoryaddrcounter_3[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => ReadMemoryState_ns(5), B => 
        un1_readmemoryaddrcounter_cry_7_S, Y => 
        readmemoryaddrcounter_3_Z(7));
    
    \mainProcess.PRDATA_8_0_iv_0_3[15]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(15), B => 
        Stamp1ShadowReg2_Z(15), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(15));
    
    \ControllUnitSubState_ns_i_a7_0_0[1]\ : CFG3
      generic map(INIT => x"13")

      port map(A => ConfigStatusReg_Z(2), B => 
        ControllUnitState_Z(2), C => ControllUnitState_Z(0), Y
         => ControllUnitSubState_ns_i_a7_0_Z(1));
    
    \ConfigStatusReg_RNO[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => sb_sb_0_STAMP_PWDATA(1), B => N_4348, C => 
        N_4340, Y => N_252_i);
    
    \CommandReg[29]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(29));
    
    \Command_RNO[4]\ : CFG2
      generic map(INIT => x"2")

      port map(A => sb_sb_0_STAMP_PWDATA(28), B => 
        SPIState_RNI27U44_Z(1), Y => N_172_i);
    
    \mainProcess.PRDATA_8_0_iv_0_1[29]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ConfigStatusReg_Z(29), B => CommandReg_Z(29), 
        C => N_1025, D => N_4335, Y => PRDATA_8_0_iv_0_1(29));
    
    \mainProcess.InternalAddr2Memory_34_1[2]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => readmemorylimitedcnt_Z(2), B => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), C => N_138, Y
         => InternalAddr2Memory_34_1(2));
    
    \CurrentAddrReg[20]\ : SLE
      port map(D => un1_currentaddrreg_cry_20_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(20));
    
    \tempcounter[7]\ : SLE
      port map(D => tempcounter_7_iv_i(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_enabletimestampgen2_1_i, ALn
         => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, 
        LAT => \GND\, Q => tempcounter_Z(7));
    
    \ControllUnitState_ns_0_0[0]\ : CFG4
      generic map(INIT => x"FF45")

      port map(A => ConfigStatusReg_Z(2), B => 
        ControllUnitState_Z(0), C => N_4344, D => 
        ControllUnitState_Z(1), Y => ControllUnitState_ns(0));
    
    \un23_0_0[2]\ : CFG4
      generic map(INIT => x"FEC0")

      port map(A => ControllUnitState_Z(3), B => 
        ControllUnitSubState_Z(1), C => N_4351, D => 
        ControllUnitSubState_Z(0), Y => un23_0_0_Z(2));
    
    \readmemoryaddrcounter[24]\ : SLE
      port map(D => readmemoryaddrcounter_3_Z(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \GND\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemoryaddrcounter_Z(24));
    
    \Stamp1ShadowReg2[24]\ : SLE
      port map(D => STAMP_0_data_frame(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(24));
    
    \ControllUnitState[10]\ : SLE
      port map(D => ControllUnitState_Z(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(10));
    
    \StartAddrReg[4]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(4));
    
    \readmemorylimitedcnt[2]\ : SLE
      port map(D => readmemorylimitedcnt_5(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorylimitedcnt_Z(2));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[6]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(6), B => TimeStampValue(6), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(6));
    
    \SPITransmitReg[10]\ : SLE
      port map(D => SPITransmitReg_13(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(10));
    
    un1_enabletimestampgen2_5_6 : CFG3
      generic map(INIT => x"C8")

      port map(A => ControllUnitState_Z(4), B => N_4343_i, C => 
        ControllUnitState_Z(7), Y => 
        un1_enabletimestampgen2_5_6_Z);
    
    un1_currentaddrreg_cry_17 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(17), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_16_Z, S => 
        un1_currentaddrreg_cry_17_S, Y => 
        un1_currentaddrreg_cry_17_Y, FCO => 
        un1_currentaddrreg_cry_17_Z);
    
    \PRDATA[1]\ : SLE
      port map(D => PRDATA_8(1), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(1));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[9]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(9), C => 
        Stamp1ShadowReg2_Z(9), D => 
        InternalData2Memory_27_0_iv_0_1(9), Y => 
        InternalData2Memory_27(9));
    
    \mainProcess.PRDATA_8_0_iv_0_0[26]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(26), D => SPIRecReg(26), Y => 
        PRDATA_8_0_iv_0_0(26));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[5]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(5), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(5));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[15]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(15), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(15));
    
    \mainProcess.PRDATA_8_0_iv_0_0[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(30), D => SPIRecReg(30), Y => 
        PRDATA_8_0_iv_0_0(30));
    
    \mainProcess.InternalAddr2Memory_34_m2[1]\ : CFG4
      generic map(INIT => x"C7C2")

      port map(A => ControllUnitState_Z(2), B => 
        InternalAddr2Memory_34_m2_1_1(1), C => 
        InternalAddr2Memory_34_sm0, D => un1_memorycnt_1_cry_1_Y, 
        Y => InternalAddr2Memory_34_m2(1));
    
    \StampFSMR1[15]\ : SLE
      port map(D => pageaddr_5_i_m4(15), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(15));
    
    \ControllUnitState_ns_0_0_o4[12]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_4342, B => N_5700, Y => N_4353);
    
    \Stamp1ShadowReg1[4]\ : SLE
      port map(D => STAMP_0_data_frame(36), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(4));
    
    \ControllUnitState_ns_0_0[8]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ControllUnitState_Z(7), B => 
        ControllUnitState_Z(6), C => N_4339, D => N_1045, Y => 
        ControllUnitState_ns(8));
    
    un1_currentaddrreg_cry_9 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(9), B => pageaddr(9), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_8_Z, S
         => un1_currentaddrreg_cry_9_S, Y => 
        un1_currentaddrreg_cry_9_Y, FCO => 
        un1_currentaddrreg_cry_9_Z);
    
    \mainProcess.pageaddr_5_i_m4[12]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(12), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(12), Y => pageaddr_5_i_m4(12));
    
    \Command[5]\ : SLE
      port map(D => N_170_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        Command_1_sqmuxa_1_i_Z, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        Command_Z(5));
    
    \readmemorycounter_RNI7QMT[1]\ : CFG2
      generic map(INIT => x"7")

      port map(A => readmemorycounter_Z(0), B => 
        readmemorycounter_Z(1), Y => N_4268);
    
    \mainProcess.InternalAddr2Memory_34_m0[6]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ControllUnitState_Z(2), B => 
        un1_memorycnt_1_cry_6_S, C => StampFSMPC_Z(6), Y => 
        InternalAddr2Memory_34_m0(6));
    
    \readmemoryaddrcounter[23]\ : SLE
      port map(D => readmemoryaddrcounter_3_Z(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemoryaddrcounter_Z(23));
    
    \Stamp1ShadowReg1[30]\ : SLE
      port map(D => STAMP_0_data_frame(62), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(30));
    
    \mainProcess.ConfigStatusReg_26_i_m2[1]\ : CFG4
      generic map(INIT => x"3AAA")

      port map(A => ConfigStatusReg_Z(1), B => SPIaddr_Z(0), C
         => ControllUnitState_Z(1), D => GPIO_6_M2F_c, Y => 
        N_4348);
    
    \ReadMemoryShadowReg[5]\ : SLE
      port map(D => InternalDataFromMem(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(5));
    
    \PRDATA[31]\ : SLE
      port map(D => PRDATA_8(31), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(31));
    
    \ConfigStatusReg_RNO_1[29]\ : CFG4
      generic map(INIT => x"F404")

      port map(A => SPIState_ns(3), B => ConfigStatusReg_Z(29), C
         => GPIO_6_M2F_c, D => m94_1_1, Y => N_149_mux);
    
    \CommandReg[19]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(19));
    
    \Stamp1ShadowReg2[2]\ : SLE
      port map(D => STAMP_0_data_frame(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(2));
    
    \mainProcess.PRDATA_8_0_iv_0_6[24]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(24), C => 
        PRDATA_8_0_iv_0_1(24), D => PRDATA_8_0_iv_0_0(24), Y => 
        PRDATA_8_0_iv_0_6(24));
    
    \ControllUnitState_ns_i_0_2[11]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => ControllUnitState_Z(4), B => 
        ConfigStatusReg_Z(2), C => 
        ControllUnitState_ns_i_0_1_Z(11), D => N_1041, Y => 
        ControllUnitState_ns_i_0_2_Z(11));
    
    \ControllUnitState_ns_i_0_a4[11]\ : CFG2
      generic map(INIT => x"1")

      port map(A => ControllUnitState_Z(3), B => 
        ControllUnitState_Z(4), Y => N_1041);
    
    un8_tempcounter_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => StampFSMPC_Z(2), C => \GND\, D
         => \GND\, FCI => un8_tempcounter_cry_1_Z, S => 
        un8_tempcounter_cry_2_S, Y => un8_tempcounter_cry_2_Y, 
        FCO => un8_tempcounter_cry_2_Z);
    
    un1_APBState_1_1_0_0_a2 : CFG3
      generic map(INIT => x"E0")

      port map(A => sb_sb_0_STAMP_PADDR(4), B => 
        sb_sb_0_STAMP_PADDR(5), C => sb_sb_0_STAMP_PADDR(6), Y
         => N_4546);
    
    \SPITransmitReg_RNO[14]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_17, B => InternalDataFromMem(14), C => 
        N_54, D => N_15_mux_16, Y => SPITransmitReg_13(14));
    
    \readmemorycounter[1]\ : SLE
      port map(D => readmemorycounter_6(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorycounter_Z(1));
    
    \mainProcess.PRDATA_8_0_iv_0_3[7]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(7), B => 
        Stamp1ShadowReg2_Z(7), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(7));
    
    \SPITransmitReg_RNO_0[31]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(23), Y => N_4_0);
    
    \PRDATA[16]\ : SLE
      port map(D => PRDATA_8(16), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(16));
    
    \InternalData2Memory[27]\ : SLE
      port map(D => InternalData2Memory_27(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(27));
    
    \SPITransmitReg_RNO_1[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_4272_i, B => ReadMemoryState_Z(8), Y => 
        SPITransmitReg_RNO_1_Z(4));
    
    \mainProcess.PRDATA_8_0_iv_0_0[3]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(3), D => SPIRecReg(3), Y => 
        PRDATA_8_0_iv_0_0(3));
    
    \StartAddrReg[14]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(14));
    
    un1_APBState_1_1_RNI4J6L : CFG4
      generic map(INIT => x"0001")

      port map(A => N_4546, B => N_4547, C => un1_APBState_1_1_Z, 
        D => un1_APBState_1_2_0_Z, Y => un1_APBState_1_i);
    
    \CurrentAddrReg[15]\ : SLE
      port map(D => un1_currentaddrreg_cry_15_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(15));
    
    \ReadMemoryState_ns_i_0_a3_2_8[3]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => ReadMemoryState_Z(6), B => 
        readmemoryaddrcounter_Z(25), C => 
        ReadMemoryState_ns_i_0_a3_2_6_Z(3), D => 
        ReadMemoryState_Z(5), Y => 
        ReadMemoryState_ns_i_0_a3_2_8_Z(3));
    
    \mainProcess.PRDATA_8_0_iv_0_2[21]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(21), 
        D => CurrentAddrReg_Z(21), Y => PRDATA_8_0_iv_0_2(21));
    
    \MemoryPageSize[3]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(3));
    
    \Stamp1ShadowReg1[6]\ : SLE
      port map(D => STAMP_0_data_frame(38), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(6));
    
    \mainProcess.PRDATA_8_0_iv_0_1[17]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ConfigStatusReg_Z(17), B => CommandReg_Z(17), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(17));
    
    \ReadMemoryState_RNO[8]\ : CFG4
      generic map(INIT => x"8ACF")

      port map(A => ReadMemoryState_Z(8), B => 
        ReadMemoryState_Z(0), C => N_2471_i_1, D => N_2496, Y => 
        N_2471_i);
    
    \ReadMemoryShadowReg[2]\ : SLE
      port map(D => InternalDataFromMem(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(2));
    
    \mainProcess.InternalAddr2Memory_34[4]\ : CFG4
      generic map(INIT => x"FDDD")

      port map(A => InternalAddr2Memory_34_1(4), B => 
        InternalAddr2Memory_34_6, C => 
        readmemoryaddrcounter_Z(27), D => ReadMemoryState_Z(4), Y
         => InternalAddr2Memory_34(4));
    
    \SPITransmitReg_RNO[1]\ : CFG4
      generic map(INIT => x"FBFA")

      port map(A => N_13_mux_0, B => N_54, C => 
        SPITransmitReg_RNO_1_Z(1), D => InternalDataFromMem(1), Y
         => SPITransmitReg_13(1));
    
    \StampFSMPC[4]\ : SLE
      port map(D => StampFSMPC_6(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_1246_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => StampFSMPC_Z(4));
    
    \mainProcess.InternalData2Memory_27_0_iv[24]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_2(24), C => 
        Stamp1ShadowReg2_Z(24), D => 
        InternalData2Memory_27_0_iv_0(24), Y => 
        InternalData2Memory_27(24));
    
    \mainProcess.PRDATA_8_0_iv_0_2[15]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(15), 
        D => CurrentAddrReg_Z(15), Y => PRDATA_8_0_iv_0_2(15));
    
    \ControllUnitState_ns_i_0_o4[14]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_4344, B => N_4342, C => dataReady_0, D => 
        ControllUnitState_Z(3), Y => N_4350);
    
    \SPITransmitReg_RNO_1[9]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(9), Y => N_15_mux_21);
    
    \SPITransmitReg[26]\ : SLE
      port map(D => SPITransmitReg_13(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(26));
    
    \CurrentAddrReg[24]\ : SLE
      port map(D => un1_currentaddrreg_cry_24_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(24));
    
    \SPITransmitReg_RNO_0[20]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(12), Y => N_4_11);
    
    \SPITransmitReg_RNO_1[18]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(18), Y => N_15_mux_12);
    
    \Command[7]\ : SLE
      port map(D => N_166_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        Command_1_sqmuxa_1_i_Z, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        Command_Z(7));
    
    \PRDATA[2]\ : SLE
      port map(D => PRDATA_8(2), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(2));
    
    \CurrentAddrReg[7]\ : SLE
      port map(D => un1_currentaddrreg_cry_7_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(7));
    
    \ControllUnitSubState_RNO[1]\ : CFG4
      generic map(INIT => x"0111")

      port map(A => N_2641, B => ControllUnitSubState_ns_i_2_Z(1), 
        C => ControllUnitSubState_ns_i_a7_4_5_Z(1), D => 
        ControllUnitSubState_ns_i_a7_4_4_Z(1), Y => N_2629_i);
    
    \StampFSMPC[5]\ : SLE
      port map(D => StampFSMPC_6(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_1246_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => StampFSMPC_Z(5));
    
    \readmemoryaddrcounter[31]\ : SLE
      port map(D => readmemoryaddrcounter_3_Z(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemoryaddrcounter_Z(31));
    
    \mainProcess.PRDATA_8_0_iv_0_2[3]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(3), 
        D => CurrentAddrReg_Z(3), Y => PRDATA_8_0_iv_0_2(3));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[28]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(28), B => 
        TimeStampValue(28), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(28));
    
    \InternalData2Memory[14]\ : SLE
      port map(D => InternalData2Memory_27(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(14));
    
    \mainProcess.PRDATA_8_0_iv_0_0[6]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(6), D => SPIRecReg(6), Y => 
        PRDATA_8_0_iv_0_0(6));
    
    \mainProcess.PRDATA_8_0_iv_0_0[28]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(28), D => SPIRecReg(28), Y => 
        PRDATA_8_0_iv_0_0(28));
    
    un1_readmemoryaddrcounter_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemoryaddrcounter_Z(28), C
         => \GND\, D => \GND\, FCI => 
        un1_readmemoryaddrcounter_cry_2_Z, S => 
        un1_readmemoryaddrcounter_cry_3_S, Y => 
        un1_readmemoryaddrcounter_cry_3_Y, FCO => 
        un1_readmemoryaddrcounter_cry_3_Z);
    
    \mainProcess.ConfigStatusReg_26_0_a2_1_RNO[30]\ : CFG4
      generic map(INIT => x"2F0F")

      port map(A => N_1316_i, B => ControllUnitState_Z(14), C => 
        GPIO_6_M2F_c, D => ConfigStatusReg_24_sn_N_5, Y => 
        ConfigStatusReg_24_sn_N_11_mux);
    
    \mainProcess.PRDATA_8_0_iv_0_1[5]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ConfigStatusReg_Z(5), B => CommandReg_Z(5), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(5));
    
    \ConfigStatusReg_RNO_0[3]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => m86_m7_0, B => r_N_6_mux, C => m84_m7_0, D
         => sb_sb_0_STAMP_PADDR(11), Y => m86_0_1);
    
    \mainProcess.PRDATA_8_0_iv_0_1[31]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ConfigStatusReg_Z(31), B => CommandReg_Z(31), 
        C => N_1025, D => N_4335, Y => PRDATA_8_0_iv_0_1(31));
    
    \ConfigStatusReg[6]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(6));
    
    ReadMemoryShadowReg_0_sqmuxa_i : CFG2
      generic map(INIT => x"E")

      port map(A => APB3ReadMemoryLimitedState_Z(3), B => 
        ReadMemoryState_Z(1), Y => 
        ReadMemoryShadowReg_0_sqmuxa_i_Z);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[20]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(20), C => pageaddr(28), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(20));
    
    \mainProcess.PRDATA_8_0_iv_0_3[10]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(10), B => 
        Stamp1ShadowReg2_Z(10), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(10));
    
    \mainProcess.PRDATA_8_0_iv_0_3[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(30), B => 
        Stamp1ShadowReg2_Z(30), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(30));
    
    \ReadMemoryShadowReg[31]\ : SLE
      port map(D => InternalDataFromMem(31), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(31));
    
    \ConfigStatusReg_RNO_3[29]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ConfigStatusReg_Z(29), B => SPIState_Z(2), C
         => counter9, Y => N_89);
    
    \mainProcess.PRDATA_8_0_iv_0_0[2]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(2), D => SPIRecReg(2), Y => 
        PRDATA_8_0_iv_0_0(2));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[19]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(19), C => 
        Stamp1ShadowReg2_Z(19), D => 
        InternalData2Memory_27_0_iv_0_1(19), Y => 
        InternalData2Memory_27(19));
    
    \StampFSMR1[26]\ : SLE
      port map(D => pageaddr_5_i_m4(26), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(26));
    
    \mainProcess.pageaddr_5_i_m4[11]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(11), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(11), Y => pageaddr_5_i_m4(11));
    
    \mainProcess.PRDATA_8_0_iv_0[20]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(20), B => 
        PRDATA_8_0_iv_0_3(20), C => PRDATA_8_0_iv_0_6(20), Y => 
        PRDATA_8(20));
    
    \mainProcess.InternalAddr2Memory_34_m2_1_0[8]\ : CFG3
      generic map(INIT => x"1B")

      port map(A => ControllUnitState_Z(2), B => 
        un1_memorycnt_1_s_8_S, C => StampFSMPC_Z(8), Y => 
        InternalAddr2Memory_34_m2_1_0(8));
    
    \readmemorycounter[0]\ : SLE
      port map(D => N_4260_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => readmemorycounter_Z(0));
    
    \ControllUnitState_ns_i_0_m2[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => ControllUnitSubState_Z(0), B => 
        ControllUnitState_Z(4), C => ControllUnitSubState_Z(1), Y
         => N_4423);
    
    \Stamp1ShadowReg1[28]\ : SLE
      port map(D => STAMP_0_data_frame(60), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(28));
    
    \mainProcess.PRDATA_8_0_iv_0_6[8]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(8), C => 
        PRDATA_8_0_iv_0_1(8), D => PRDATA_8_0_iv_0_0(8), Y => 
        PRDATA_8_0_iv_0_6(8));
    
    \mainProcess.InternalData2Memory_27_0_iv_3[11]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(11), B => 
        TimeStampValue(11), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_3(11));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(1), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(1));
    
    un1_currentaddrreg_cry_28 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(28), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_27_Z, S => 
        un1_currentaddrreg_cry_28_S, Y => 
        un1_currentaddrreg_cry_28_Y, FCO => 
        un1_currentaddrreg_cry_28_Z);
    
    \mainProcess.PRDATA_8_0_iv_0_1[2]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ConfigStatusReg_Z(2), B => CommandReg_Z(2), C
         => N_1025, D => N_4335, Y => PRDATA_8_0_iv_0_1(2));
    
    \mainProcess.PRDATA_8_0_iv_0[2]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(2), B => 
        PRDATA_8_0_iv_0_3(2), C => PRDATA_8_0_iv_0_6(2), Y => 
        PRDATA_8(2));
    
    \mainProcess.PRDATA_8_0_iv_0_6[7]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(7), C => 
        PRDATA_8_0_iv_0_1(7), D => PRDATA_8_0_iv_0_0(7), Y => 
        PRDATA_8_0_iv_0_6(7));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[14]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(14), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(14));
    
    \InternalData2Memory[1]\ : SLE
      port map(D => InternalData2Memory_27(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(1));
    
    \Command[0]\ : SLE
      port map(D => N_180_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        Command_1_sqmuxa_1_i_Z, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        Command_Z(0));
    
    un1_readmemoryaddrcounter_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemoryaddrcounter_Z(25), C
         => \GND\, D => \GND\, FCI => 
        un1_readmemoryaddrcounter_cry_5_Z, S => 
        un1_readmemoryaddrcounter_cry_6_S, Y => 
        un1_readmemoryaddrcounter_cry_6_Y, FCO => 
        un1_readmemoryaddrcounter_cry_6_Z);
    
    \ControllUnitState_ns_i_a2_1[11]\ : CFG2
      generic map(INIT => x"1")

      port map(A => memorycnt_Z(1), B => memorycnt_Z(2), Y => 
        N_2624_1);
    
    \ConfigStatusReg_RNO_0[2]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => m87_m7_0, B => r_N_6_mux, C => m84_m7_0, D
         => sb_sb_0_STAMP_PADDR(11), Y => m87_0_1);
    
    \SPITransmitReg[2]\ : SLE
      port map(D => SPITransmitReg_13(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(2));
    
    \ReadMemoryShadowReg[13]\ : SLE
      port map(D => InternalDataFromMem(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(13));
    
    \mainProcess.PRDATA_8_0_iv_0_3[12]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(12), B => 
        Stamp1ShadowReg2_Z(12), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(12));
    
    \CurrentAddrReg[26]\ : SLE
      port map(D => un1_currentaddrreg_cry_26_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(26));
    
    \CurrentAddrReg[2]\ : SLE
      port map(D => un1_currentaddrreg_cry_2_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(2));
    
    \isfirstrun_RNO[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => ControllUnitState_RNI2VHT_Z(14), B => 
        isfirstrun_Z(0), Y => isfirstrun_1_sqmuxa);
    
    \APB3ReadMemoryLimitedState[2]\ : SLE
      port map(D => N_101, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => APB3ReadMemoryLimitedState_Z(2));
    
    \MemoryPageSize[8]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(8));
    
    \mainProcess.InternalAddr2Memory_34[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => InternalAddr2Memory_34_m5(0), B => N_143_mux, 
        C => InternalAddr2Memory_34_m2(0), Y => 
        InternalAddr2Memory_34(0));
    
    enableTimestampGen : SLE
      port map(D => GPIO_6_M2F_c, CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => enableTimestampGen_Z);
    
    \MemoryPageSize[5]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(5));
    
    \mainProcess.PRDATA_8_0_iv_0_3[13]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(13), B => 
        Stamp1ShadowReg2_Z(13), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(13));
    
    SPIaddr_2_sqmuxa_1_i_m2 : CFG4
      generic map(INIT => x"C5F5")

      port map(A => ControllUnitState_Z(1), B => isfirstrun_Z(0), 
        C => ControllUnitState_Z(14), D => dataReady_0, Y => 
        N_4424);
    
    \SPITransmitReg_RNO_1[30]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(30), Y => N_15_mux_0);
    
    \mainProcess.PRDATA_8_0_iv_0_a2_11[12]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => sb_sb_0_STAMP_PADDR(3), B => 
        sb_sb_0_STAMP_PADDR(4), C => sb_sb_0_STAMP_PADDR(6), D
         => sb_sb_0_STAMP_PADDR(5), Y => N_1033);
    
    \mainProcess.InternalAddr2Memory_34_m2[0]\ : CFG3
      generic map(INIT => x"AB")

      port map(A => ControllUnitState_Z(11), B => 
        InternalAddr2Memory_34_m2_1_1(0), C => 
        InternalAddr2Memory_34_sm0, Y => 
        InternalAddr2Memory_34_m2(0));
    
    \mainProcess.pageaddr_5_i_m4[9]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(9), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(9), Y => pageaddr_5_i_m4(9));
    
    \StampFSMR1[25]\ : SLE
      port map(D => pageaddr_5_i_m4(25), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(25));
    
    \ReadMemoryState_ns_i_0_a3_2_6[3]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => readmemoryaddrcounter_Z(30), B => 
        readmemoryaddrcounter_Z(27), C => 
        readmemoryaddrcounter_Z(24), D => 
        readmemoryaddrcounter_Z(23), Y => 
        ReadMemoryState_ns_i_0_a3_2_6_Z(3));
    
    \mainProcess.PRDATA_8_0_iv_0[31]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(31), B => 
        PRDATA_8_0_iv_0_3(31), C => PRDATA_8_0_iv_0_6(31), Y => 
        PRDATA_8(31));
    
    \mainProcess.InternalAddr2Memory_34_m5[0]\ : CFG4
      generic map(INIT => x"880F")

      port map(A => readmemorylimitedcnt_Z(0), B => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), C => N_4258, D
         => N_138, Y => InternalAddr2Memory_34_m5(0));
    
    \memorycnt[3]\ : SLE
      port map(D => memorycnt_6(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => memorycnt_Z(3));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[26]\ : CFG4
      generic map(INIT => x"ACA0")

      port map(A => SPIRecReg(26), B => pageaddr(2), C => 
        ReadMemoryState_Z(4), D => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0(26));
    
    \tempcounter[3]\ : SLE
      port map(D => N_4295_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_enabletimestampgen2_1_i, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tempcounter_Z(3));
    
    \ReadMemoryState_ns_0_a3_0_a3[5]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => readmemoryaddrcounter_Z(25), B => 
        ReadMemoryState_ns_i_0_a3_2_6_Z(3), C => 
        ReadMemoryState_ns_i_0_a3_2_7_Z(3), D => 
        ReadMemoryState_Z(4), Y => ReadMemoryState_ns(5));
    
    \ReadMemoryShadowReg[30]\ : SLE
      port map(D => InternalDataFromMem(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(30));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[27]\ : CFG4
      generic map(INIT => x"ACA0")

      port map(A => SPIRecReg(27), B => pageaddr(3), C => 
        ReadMemoryState_Z(4), D => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0(27));
    
    \Stamp1ShadowReg1[12]\ : SLE
      port map(D => STAMP_0_data_frame(44), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(12));
    
    \InternalData2Memory[12]\ : SLE
      port map(D => InternalData2Memory_27(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(12));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[10]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(10), C => pageaddr(18), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(10));
    
    \SPITransmitReg[4]\ : SLE
      port map(D => SPITransmitReg_13(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(4));
    
    \mainProcess.pageaddr_5_i_m4[23]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(23), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(23), Y => pageaddr_5_i_m4(23));
    
    \ReadMemoryShadowReg[25]\ : SLE
      port map(D => InternalDataFromMem(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(25));
    
    \mainProcess.PRDATA_8_0_iv_0_0[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(4), D => SPIRecReg(4), Y => 
        PRDATA_8_0_iv_0_0(4));
    
    \ReadMemoryShadowReg[3]\ : SLE
      port map(D => InternalDataFromMem(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(3));
    
    \mainProcess.PRDATA_8_0_iv_0_1[26]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ConfigStatusReg_Z(26), B => CommandReg_Z(26), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(26));
    
    \mainProcess.InternalData2Memory_27_0_iv_2[30]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(30), B => 
        TimeStampValue(30), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_2(30));
    
    ControllUnitState_8_sqmuxa_i_o3_0 : CFG2
      generic map(INIT => x"7")

      port map(A => GPIO_6_M2F_c, B => ControllUnitSubState_Z(1), 
        Y => N_1257_i);
    
    \mainProcess.PRDATA_8_0_iv_0[16]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(16), B => 
        PRDATA_8_0_iv_0_3(16), C => PRDATA_8_0_iv_0_6(16), Y => 
        PRDATA_8(16));
    
    \APBState_RNIE91K[1]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => sb_sb_0_STAMP_PADDR(7), B => 
        sb_sb_0_STAMP_PADDR(10), C => APBState_Z(1), D => 
        sb_sb_0_STAMP_PADDR(11), Y => SPIState_m2_e_1);
    
    \mainProcess.PRDATA_8_0_iv_0_3[25]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(25), B => 
        Stamp1ShadowReg2_Z(25), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(25));
    
    Command_1_sqmuxa_0_a2_1 : CFG3
      generic map(INIT => x"10")

      port map(A => un1_APBState_1_2_0_Z, B => 
        sb_sb_0_STAMP_PADDR(11), C => Command_1_sqmuxa_0_a2_1_0_Z, 
        Y => N_1186);
    
    \APBState_ns_1_0_.m5_0_a2\ : CFG4
      generic map(INIT => x"0800")

      port map(A => sb_sb_0_STAMP_PENABLE, B => 
        sb_sb_0_Memory_PSELx, C => N_1539_i, D => 
        sb_sb_0_STAMP_PWRITE, Y => APBState_ns(1));
    
    \mainProcess.InternalAddr2Memory_34[3]\ : CFG4
      generic map(INIT => x"FDDD")

      port map(A => InternalAddr2Memory_34_1(3), B => 
        InternalAddr2Memory_34_14, C => 
        readmemoryaddrcounter_Z(28), D => ReadMemoryState_Z(4), Y
         => InternalAddr2Memory_34(3));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[8]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(8), B => TimeStampValue(8), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(8));
    
    \mainProcess.PRDATA_8_0_iv_0_0[21]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(21), D => SPIRecReg(21), Y => 
        PRDATA_8_0_iv_0_0(21));
    
    \mainProcess.memorycnt_6_cry_4\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => N_1541_i, C => memorycnt_Z(5), D
         => \GND\, FCI => memorycnt_6_cry_3, S => memorycnt_6(5), 
        Y => memorycnt_6_cry_4_Y, FCO => memorycnt_6_cry_4);
    
    \mainProcess.ConfigStatusReg_26_i_o4[31]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => sb_sb_0_STAMP_PADDR(2), B => 
        sb_sb_0_STAMP_PADDR(6), C => sb_sb_0_STAMP_PADDR(3), Y
         => N_4335);
    
    \StampFSMPC_RNO[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => ControllUnitState_Z(11), B => StampFSMPC_Z(0), 
        Y => N_746_i);
    
    \SPITransmitReg_RNO[15]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_16, B => InternalDataFromMem(15), C => 
        N_54, D => N_15_mux_15, Y => SPITransmitReg_13(15));
    
    \SPITransmitReg[15]\ : SLE
      port map(D => SPITransmitReg_13(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(15));
    
    \mainProcess.memorycnt_6_cry_2_0\ : ARI1
      generic map(INIT => x"52122")

      port map(A => ControllUnitState_Z(3), B => memorycnt_Z(3), 
        C => ControllUnitState_RNI2VHT_Z(14), D => N_1255_i, FCI
         => memorycnt_6_cry_1, S => memorycnt_6(3), Y => 
        memorycnt_6_cry_2_0_Y, FCO => memorycnt_6_cry_2);
    
    \memorycnt[5]\ : SLE
      port map(D => memorycnt_6(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => memorycnt_Z(5));
    
    un1_readmemoryaddrcounter_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemoryaddrcounter_Z(29), C
         => \GND\, D => \GND\, FCI => 
        un1_readmemoryaddrcounter_cry_1_Z, S => 
        un1_readmemoryaddrcounter_cry_2_S, Y => 
        un1_readmemoryaddrcounter_cry_2_Y, FCO => 
        un1_readmemoryaddrcounter_cry_2_Z);
    
    \SPITransmitReg_RNO_0[1]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(1), Y => N_13_mux_0);
    
    SPITransmitReg_0_sqmuxa_2_i_m2 : CFG4
      generic map(INIT => x"CCC5")

      port map(A => ReadMemoryState_Z(6), B => N_4272_i, C => 
        ReadMemoryState_Z(7), D => ReadMemoryState_Z(8), Y => 
        N_4270);
    
    \CommandReg[0]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(0));
    
    \StartAddrReg[27]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(27));
    
    \mainProcess.PRDATA_8_0_iv_0_2[10]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(10), 
        D => CurrentAddrReg_Z(10), Y => PRDATA_8_0_iv_0_2(10));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[15]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(15), C => pageaddr(23), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(15));
    
    \StartAddrReg[12]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(12));
    
    \StampFSMPC[1]\ : SLE
      port map(D => StampFSMPC_6_Z(1), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_1246_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => StampFSMPC_Z(1));
    
    \mainProcess.PRDATA_8_0_iv_0[19]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(19), B => 
        PRDATA_8_0_iv_0_3(19), C => PRDATA_8_0_iv_0_6(19), Y => 
        PRDATA_8(19));
    
    Command_1_sqmuxa_1_i_RNO_0 : CFG3
      generic map(INIT => x"04")

      port map(A => sb_sb_0_STAMP_PADDR(10), B => m73_m2_e_0_0, C
         => sb_sb_0_STAMP_PADDR(7), Y => m73_m2_e_1);
    
    \readmemorylimitedcnt_RNIBBFG2[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemorylimitedcnt_Z(4), C => 
        \GND\, D => \GND\, FCI => un1_readmemorylimitedcnt_cry_3, 
        S => readmemorylimitedcnt_RNIBBFG2_S(4), Y => 
        readmemorylimitedcnt_RNIBBFG2_Y(4), FCO => 
        un1_readmemorylimitedcnt_cry_4);
    
    \CurrentAddrReg[21]\ : SLE
      port map(D => un1_currentaddrreg_cry_21_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(21));
    
    \counter_RNO[1]\ : CFG3
      generic map(INIT => x"E6")

      port map(A => SPIState_Z(2), B => counter_Z(1), C => 
        InternalBusy, Y => N_4253_i);
    
    PRDATA_17_sqmuxa_8_RNIDUVO : CFG4
      generic map(INIT => x"0010")

      port map(A => sb_sb_0_STAMP_PADDR(9), B => 
        sb_sb_0_STAMP_PADDR(8), C => PRDATA_17_sqmuxa_8_Z, D => 
        N_4335, Y => r_N_6_mux);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[18]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(18), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(18));
    
    \PRDATA[17]\ : SLE
      port map(D => PRDATA_8(17), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(17));
    
    \mainProcess.pageaddr_5_i_m4[18]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(18), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(18), Y => N_4370);
    
    \CommandReg[23]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(23));
    
    \SPIState_RNO[4]\ : CFG4
      generic map(INIT => x"EAAA")

      port map(A => m46_1_1_0, B => SPIState_1_sqmuxa, C => m46_0, 
        D => m46_1_1, Y => N_157_mux);
    
    \APBState[1]\ : SLE
      port map(D => APBState_ns(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => APBState_Z(1));
    
    un1_memorycnt_1_cry_3 : ARI1
      generic map(INIT => x"5A9AA")

      port map(A => N_4343, B => memorycnt_Z(3), C => N_761, D
         => N_762, FCI => un1_memorycnt_1_cry_2_Z, S => 
        un1_memorycnt_1_cry_3_S, Y => un1_memorycnt_1_cry_3_Y, 
        FCO => un1_memorycnt_1_cry_3_Z);
    
    \un23_0_o4[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => ControllUnitState_Z(5), B => 
        ControllUnitState_Z(7), Y => N_4351);
    
    \SPITransmitReg_RNO_1[10]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(10), Y => N_15_mux_20);
    
    \PRDATA[18]\ : SLE
      port map(D => PRDATA_8(18), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(18));
    
    \mainProcess.PRDATA_8_0_iv_0_2[12]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(12), 
        D => CurrentAddrReg_Z(12), Y => PRDATA_8_0_iv_0_2(12));
    
    ControllUnitState_tr25_0_a2_4 : CFG3
      generic map(INIT => x"01")

      port map(A => tempcounter_Z(8), B => tempcounter_Z(5), C
         => tempcounter_Z(4), Y => 
        ControllUnitState_tr25_0_a2_4_Z);
    
    \StartAddrReg[13]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(13));
    
    \SPITransmitReg[29]\ : SLE
      port map(D => SPITransmitReg_13(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(29));
    
    \ReadMemoryState_ns_i_m3_i_o2[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => N_4272_i, B => InternalBusy, Y => N_68);
    
    \tempcounter[8]\ : SLE
      port map(D => N_4299_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_enabletimestampgen2_1_i, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tempcounter_Z(8));
    
    \readmemorycounter_RNO[2]\ : CFG4
      generic map(INIT => x"E02C")

      port map(A => N_1508_i, B => un1_enableSPI_1_sqmuxa_1_i, C
         => readmemorycounter_Z(2), D => N_4268, Y => N_4261_i);
    
    \mainProcess.InternalData2Memory_27_0_iv[25]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_3(25), C => 
        Stamp1ShadowReg2_Z(25), D => 
        InternalData2Memory_27_0_iv_1(25), Y => 
        InternalData2Memory_27(25));
    
    \mainProcess.PRDATA_8_0_iv_0_3[14]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(14), B => 
        Stamp1ShadowReg2_Z(14), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(14));
    
    \mainProcess.PRDATA_8_0_iv_0_2[13]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(13), 
        D => CurrentAddrReg_Z(13), Y => PRDATA_8_0_iv_0_2(13));
    
    \Stamp1ShadowReg2[28]\ : SLE
      port map(D => STAMP_0_data_frame(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(28));
    
    \readmemorylimitedcnt_RNIMSQE3[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemorylimitedcnt_Z(6), C => 
        \GND\, D => \GND\, FCI => un1_readmemorylimitedcnt_cry_5, 
        S => readmemorylimitedcnt_RNIMSQE3_S(6), Y => 
        readmemorylimitedcnt_RNIMSQE3_Y(6), FCO => 
        un1_readmemorylimitedcnt_cry_6);
    
    \readmemorylimitedcnt[4]\ : SLE
      port map(D => readmemorylimitedcnt_5(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorylimitedcnt_Z(4));
    
    \mainProcess.InternalData2Memory_27_0_iv[21]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_3(21), C => 
        Stamp1ShadowReg2_Z(21), D => 
        InternalData2Memory_27_0_iv_1(21), Y => 
        InternalData2Memory_27(21));
    
    \SPITransmitReg_RNO[4]\ : CFG4
      generic map(INIT => x"FBFA")

      port map(A => N_13_mux, B => N_54, C => 
        SPITransmitReg_RNO_1_Z(4), D => InternalDataFromMem(4), Y
         => SPITransmitReg_13(4));
    
    \CurrentAddrReg[27]\ : SLE
      port map(D => un1_currentaddrreg_cry_27_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(27));
    
    \StampFSMR1[19]\ : SLE
      port map(D => N_4369, CLK => sb_sb_0_FIC_0_CLK, EN => 
        ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        pageaddr(19));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[19]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(19), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(19));
    
    un1_APBState_1_5_RNIEAJU1 : CFG4
      generic map(INIT => x"0400")

      port map(A => SPIState_m2_e_1_0_Z, B => SPIState_m2_e_1, C
         => \un1_APBState_1_5_1z\, D => SPIState_m2_e_1_1_Z, Y
         => SPIState_1_sqmuxa);
    
    \mainProcess.PRDATA_8_0_iv_0_6[9]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(9), C => 
        PRDATA_8_0_iv_0_1(9), D => PRDATA_8_0_iv_0_0(9), Y => 
        PRDATA_8_0_iv_0_6(9));
    
    \SPITransmitReg_RNO_0[24]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(16), Y => N_4_7);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[1]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(1), C => pageaddr(9), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(1));
    
    \readmemorylimitedcnt[5]\ : SLE
      port map(D => readmemorylimitedcnt_5(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorylimitedcnt_Z(5));
    
    \mainProcess.PRDATA_8_0_iv_0[28]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(28), B => 
        PRDATA_8_0_iv_0_3(28), C => PRDATA_8_0_iv_0_6(28), Y => 
        PRDATA_8(28));
    
    ControllUnitSubState_2_sqmuxa_i_o3_RNIDUPQ : CFG3
      generic map(INIT => x"B0")

      port map(A => ControllUnitState_Z(11), B => N_1261_i, C => 
        GPIO_6_M2F_c, Y => N_1246_i);
    
    \StampFSMPC[8]\ : SLE
      port map(D => StampFSMPC_6(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_1246_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => StampFSMPC_Z(8));
    
    \mainProcess.PRDATA_8_0_iv_0_0[17]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(17), D => SPIRecReg(17), Y => 
        PRDATA_8_0_iv_0_0(17));
    
    \StampFSMR1[12]\ : SLE
      port map(D => pageaddr_5_i_m4(12), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(12));
    
    \Stamp1ShadowReg1[15]\ : SLE
      port map(D => STAMP_0_data_frame(47), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(15));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[0]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(0), B => TimeStampValue(0), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(0));
    
    \readmemorylimitedcnt[6]\ : SLE
      port map(D => readmemorylimitedcnt_5(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorylimitedcnt_Z(6));
    
    \mainProcess.PRDATA_8_0_iv_0_1[28]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ConfigStatusReg_Z(28), B => CommandReg_Z(28), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(28));
    
    un1_currentaddrreg_cry_6 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(6), B => pageaddr(6), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_5_Z, S
         => un1_currentaddrreg_cry_6_S, Y => 
        un1_currentaddrreg_cry_6_Y, FCO => 
        un1_currentaddrreg_cry_6_Z);
    
    \CommandReg[13]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(13));
    
    \SPITransmitReg[17]\ : SLE
      port map(D => SPITransmitReg_13(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(17));
    
    \mainProcess.PRDATA_8_0_iv_0_6[1]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(1), C => 
        PRDATA_8_0_iv_0_1(1), D => PRDATA_8_0_iv_0_0(1), Y => 
        PRDATA_8_0_iv_0_6(1));
    
    \SPITransmitReg_RNO_1[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_4272_i, B => ReadMemoryState_Z(8), Y => 
        SPITransmitReg_RNO_1_Z(1));
    
    \SPITransmitReg_RNO_1[28]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(28), Y => N_15_mux_2);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[7]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(7), B => TimeStampValue(7), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(7));
    
    \mainProcess.PRDATA_8_0_iv_0_1[15]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(7), B => CommandReg_Z(15), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(15));
    
    \CurrentAddrReg[8]\ : SLE
      port map(D => un1_currentaddrreg_cry_8_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(8));
    
    \Stamp1ShadowReg1[19]\ : SLE
      port map(D => STAMP_0_data_frame(51), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(19));
    
    \mainProcess.PRDATA_8_0_iv_0_6[17]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(17), C => 
        PRDATA_8_0_iv_0_1(17), D => PRDATA_8_0_iv_0_0(17), Y => 
        PRDATA_8_0_iv_0_6(17));
    
    \readmemoryaddrcounter_3[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => ReadMemoryState_ns(5), B => 
        un1_readmemoryaddrcounter_cry_0_S, Y => 
        readmemoryaddrcounter_3_Z(0));
    
    Command_1_sqmuxa_0_a2_1_0 : CFG2
      generic map(INIT => x"4")

      port map(A => \un1_APBState_1_5_1z\, B => APBState_Z(1), Y
         => Command_1_sqmuxa_0_a2_1_0_Z);
    
    \ReadMemoryState[1]\ : SLE
      port map(D => ReadMemoryState_Z(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ReadMemoryState_Z(1));
    
    \StartAddrReg[25]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(25));
    
    \Stamp1ShadowReg1[2]\ : SLE
      port map(D => STAMP_0_data_frame(34), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(2));
    
    \mainProcess.PRDATA_8_0_iv_0_6[29]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(29), C => 
        PRDATA_8_0_iv_0_1(29), D => PRDATA_8_0_iv_0_0(29), Y => 
        PRDATA_8_0_iv_0_6(29));
    
    \Stamp1ShadowReg2[12]\ : SLE
      port map(D => STAMP_0_data_frame(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(12));
    
    \mainProcess.PRDATA_8_0_iv_0_3[1]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(1), B => 
        Stamp1ShadowReg2_Z(1), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(1));
    
    \SPITransmitReg_RNO_0[27]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(19), Y => N_4_4);
    
    \SPITransmitReg_RNO_0[18]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(10), Y => N_4_13);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_2[31]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(31), B => 
        TimeStampValue(31), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_2(31));
    
    \mainProcess.pageaddr_5_i_m4[29]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(29), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(29), Y => pageaddr_5_i_m4(29));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[1]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(1), B => TimeStampValue(1), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(1));
    
    \CommandReg[27]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(27));
    
    \SPITransmitReg_RNO[19]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_12, B => InternalDataFromMem(19), C => 
        N_54, D => N_15_mux_11, Y => SPITransmitReg_13(19));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[29]\ : CFG4
      generic map(INIT => x"ACA0")

      port map(A => SPIRecReg(29), B => pageaddr(5), C => 
        ReadMemoryState_Z(4), D => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0(29));
    
    \ConfigStatusReg[0]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(0));
    
    \mainProcess.pageaddr_5_i_m4[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(1), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(1), Y => pageaddr_5_i_m4(1));
    
    \mainProcess.pageaddr_5_i_m4[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(5), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(5), Y => pageaddr_5_i_m4(5));
    
    \SPITransmitReg[11]\ : SLE
      port map(D => SPITransmitReg_13(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(11));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[5]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(5), C => pageaddr(13), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(5));
    
    \StampFSMPC[3]\ : SLE
      port map(D => StampFSMPC_6(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_1246_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => StampFSMPC_Z(3));
    
    \mainProcess.PRDATA_8_0_iv_0_3[20]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(20), B => 
        Stamp1ShadowReg2_Z(20), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(20));
    
    \mainProcess.PRDATA_8_0_iv_0_2[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(30), 
        D => CurrentAddrReg_Z(30), Y => PRDATA_8_0_iv_0_2(30));
    
    \counter[1]\ : SLE
      port map(D => N_4253_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        counter_Z(0), ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => counter_Z(1));
    
    \ReadMemoryShadowReg[6]\ : SLE
      port map(D => InternalDataFromMem(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(6));
    
    \ReadMemoryShadowReg[11]\ : SLE
      port map(D => InternalDataFromMem(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(11));
    
    \ControllUnitState_RNIR5I[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => ControllUnitState_Z(2), B => 
        ControllUnitState_Z(1), Y => ConfigStatusReg_24_sn_N_5);
    
    \InternalData2Memory[19]\ : SLE
      port map(D => InternalData2Memory_27(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(19));
    
    \InternalData2Memory[16]\ : SLE
      port map(D => InternalData2Memory_27(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(16));
    
    \readmemorylimitedcnt_RNITM0U3[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemorylimitedcnt_Z(7), C => 
        \GND\, D => \GND\, FCI => un1_readmemorylimitedcnt_cry_6, 
        S => readmemorylimitedcnt_RNITM0U3_S(7), Y => 
        readmemorylimitedcnt_RNITM0U3_Y(7), FCO => 
        un1_readmemorylimitedcnt_cry_7);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[14]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(14), C => pageaddr(22), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(14));
    
    \counter_RNO[0]\ : CFG4
      generic map(INIT => x"D5AA")

      port map(A => counter_Z(0), B => counter_Z(1), C => 
        InternalBusy, D => SPIState_Z(2), Y => N_140_mux_i);
    
    \mainProcess.PRDATA_8_0_iv_0[5]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(5), B => 
        PRDATA_8_0_iv_0_3(5), C => PRDATA_8_0_iv_0_6(5), Y => 
        PRDATA_8(5));
    
    \CurrentAddrReg[19]\ : SLE
      port map(D => un1_currentaddrreg_cry_19_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(19));
    
    \SPITransmitReg_RNO[13]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_18, B => InternalDataFromMem(13), C => 
        N_54, D => N_15_mux_17, Y => SPITransmitReg_13(13));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[23]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg2_Z(23), B => 
        Stamp1ShadowReg1_Z(23), C => 
        InternalData2Memory_5_sqmuxa_Z, D => 
        InternalData2Memory_4_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_1(23));
    
    \StampFSMPC_6_0_a2[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => un8_tempcounter_cry_3_S, B => 
        ControllUnitState_Z(11), Y => StampFSMPC_6(3));
    
    \CommandReg[2]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(2));
    
    \StampFSMPC[6]\ : SLE
      port map(D => StampFSMPC_6(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_1246_i, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => StampFSMPC_Z(6));
    
    \mainProcess.PRDATA_8_0_iv_0_3[22]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(22), B => 
        Stamp1ShadowReg2_Z(22), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(22));
    
    \SPIState[2]\ : SLE
      port map(D => N_42_0, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => SPIState_Z(2));
    
    \mainProcess.PRDATA_8_0_iv_0_2[14]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(14), 
        D => CurrentAddrReg_Z(14), Y => PRDATA_8_0_iv_0_2(14));
    
    \mainProcess.SPITransmitReg_13_0_iv_0[6]\ : CFG4
      generic map(INIT => x"A808")

      port map(A => N_4270, B => InternalDataFromMem(6), C => 
        SPIState_1_sqmuxa, D => sb_sb_0_STAMP_PWDATA(6), Y => 
        SPITransmitReg_13(6));
    
    \ConfigStatusReg_RNO[2]\ : CFG4
      generic map(INIT => x"5B54")

      port map(A => ReadMemoryState_Z(3), B => 
        ConfigStatusReg_Z(2), C => N_2496_i, D => m87_0_1, Y => 
        N_88);
    
    un1_APBState_1_5 : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PADDR(0), B => 
        sb_sb_0_STAMP_PADDR(1), Y => \un1_APBState_1_5_1z\);
    
    \mainProcess.PRDATA_8_0_iv_0_6[4]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(4), C => 
        PRDATA_8_0_iv_0_1(4), D => PRDATA_8_0_iv_0_0(4), Y => 
        PRDATA_8_0_iv_0_6(4));
    
    \readmemorylimitedcnt[8]\ : SLE
      port map(D => readmemorylimitedcnt_5(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorylimitedcnt_Z(8));
    
    MemoryPageSize_1_sqmuxa_0_o4_0_RNIPMOK : CFG4
      generic map(INIT => x"0002")

      port map(A => PRDATA_17_sqmuxa_8_Z, B => 
        un1_APBState_1_2_0_Z, C => sb_sb_0_STAMP_PADDR(11), D => 
        MemoryPageSize_1_sqmuxa_0_o4_0_Z, Y => N_4340_i);
    
    un1_currentaddrreg_cry_18 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(18), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_17_Z, S => 
        un1_currentaddrreg_cry_18_S, Y => 
        un1_currentaddrreg_cry_18_Y, FCO => 
        un1_currentaddrreg_cry_18_Z);
    
    \memorycnt[7]\ : SLE
      port map(D => memorycnt_6(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => N_2624_2);
    
    \SPIState[3]\ : SLE
      port map(D => N_70, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => SPIState_Z(3));
    
    \mainProcess.pageaddr_5_i_m4[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(7), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(7), Y => pageaddr_5_i_m4(7));
    
    \SPITransmitReg_RNO[20]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_11, B => InternalDataFromMem(20), C => 
        N_54, D => N_15_mux_10, Y => SPITransmitReg_13(20));
    
    \SPITransmitReg_RNO_0[26]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(18), Y => N_4_5);
    
    \mainProcess.PRDATA_8_0_iv_0_3[23]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(23), B => 
        Stamp1ShadowReg2_Z(23), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(23));
    
    \Command_RNO[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => SPIState_RNI27U44_Z(1), B => 
        sb_sb_0_STAMP_PWDATA(25), Y => N_178_i);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[28]\ : CFG4
      generic map(INIT => x"FDEC")

      port map(A => ReadMemoryState_Z(4), B => N_4535, C => 
        SPIRecReg(28), D => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(28));
    
    \CommandReg[17]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(17));
    
    \mainProcess.PRDATA_8_0_iv_0_1[6]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ConfigStatusReg_Z(6), B => CommandReg_Z(6), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(6));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[5]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(5), C => 
        Stamp1ShadowReg2_Z(5), D => 
        InternalData2Memory_27_0_iv_0_1(5), Y => 
        InternalData2Memory_27(5));
    
    \ConfigStatusReg[23]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize(15));
    
    \mainProcess.InternalData2Memory_27_0_iv[26]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_2(26), C => 
        Stamp1ShadowReg2_Z(26), D => 
        InternalData2Memory_27_0_iv_0(26), Y => 
        InternalData2Memory_27(26));
    
    \mainProcess.PRDATA_8_0_iv_0_0[7]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(7), D => SPIRecReg(7), Y => 
        PRDATA_8_0_iv_0_0(7));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[9]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(9), C => pageaddr(17), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(9));
    
    \CurrentAddrReg[6]\ : SLE
      port map(D => un1_currentaddrreg_cry_6_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(6));
    
    \CommandReg[8]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(8));
    
    \mainProcess.PRDATA_8_0_iv_0_1[21]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(13), B => CommandReg_Z(21), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(21));
    
    \ConfigStatusReg_RNO_4[29]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_4343_i, B => ControllUnitState_Z(2), Y => 
        N_146);
    
    \Command_RNI6AH02[1]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => Command_Z(1), B => m17_e_1, C => Command_Z(3), 
        D => Command_Z(2), Y => N_21_0);
    
    \StartAddrReg[5]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(5));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[2]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(2), B => TimeStampValue(2), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(2));
    
    \ReadMemoryShadowReg[8]\ : SLE
      port map(D => InternalDataFromMem(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(8));
    
    \ReadMemoryShadowReg[10]\ : SLE
      port map(D => InternalDataFromMem(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(10));
    
    \ControllUnitSubState_ns_i_2[1]\ : CFG4
      generic map(INIT => x"F0F8")

      port map(A => N_2648, B => 
        ControllUnitSubState_ns_i_a7_0_Z(1), C => 
        ControllUnitSubState_ns_i_1_Z(1), D => N_2631, Y => 
        ControllUnitSubState_ns_i_2_Z(1));
    
    \ControllUnitState_ns_0_0[9]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ControllUnitState_Z(6), B => 
        ControllUnitState_Z(5), C => N_1045, D => N_4339, Y => 
        ControllUnitState_ns(9));
    
    \ConfigStatusReg[29]\ : SLE
      port map(D => ConfigStatusReg_40(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ConfigStatusReg_Z(29));
    
    un1_memorycnt_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => N_2624_2, C => \GND\, D => \GND\, 
        FCI => un1_memorycnt_1_cry_6_Z, S => 
        un1_memorycnt_1_cry_7_S, Y => un1_memorycnt_1_cry_7_Y, 
        FCO => un1_memorycnt_1_cry_7_Z);
    
    \mainProcess.readmemorylimitedcnt_5[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => readmemorylimitedcnt_RNI7K912_S(3), B => 
        APB3ReadMemoryLimitedState_Z(1), Y => 
        readmemorylimitedcnt_5(3));
    
    \CommandReg[22]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(22));
    
    un1_memorycnt_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => memorycnt_Z(5), C => \GND\, D => 
        \GND\, FCI => un1_memorycnt_1_cry_4_Z, S => 
        un1_memorycnt_1_cry_5_S, Y => un1_memorycnt_1_cry_5_Y, 
        FCO => un1_memorycnt_1_cry_5_Z);
    
    \InternalAddr2Memory[6]\ : SLE
      port map(D => InternalAddr2Memory_34(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => InternalAddr2Memory_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => InternalAddr2Memory_Z(6));
    
    \ConfigStatusReg_RNO_1[2]\ : CFG4
      generic map(INIT => x"0110")

      port map(A => sb_sb_0_STAMP_PADDR(7), B => 
        sb_sb_0_STAMP_PADDR(10), C => ConfigStatusReg_Z(2), D => 
        sb_sb_0_STAMP_PWDATA(2), Y => m87_m7_0);
    
    un1_currentaddrreg_cry_26 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(26), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_25_Z, S => 
        un1_currentaddrreg_cry_26_S, Y => 
        un1_currentaddrreg_cry_26_Y, FCO => 
        un1_currentaddrreg_cry_26_Z);
    
    \mainProcess.PRDATA_8_0_iv_0[14]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(14), B => 
        PRDATA_8_0_iv_0_3(14), C => PRDATA_8_0_iv_0_6(14), Y => 
        PRDATA_8(14));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[14]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(14), C => 
        Stamp1ShadowReg2_Z(14), D => 
        InternalData2Memory_27_0_iv_0_1(14), Y => 
        InternalData2Memory_27(14));
    
    \ConfigStatusReg[25]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(25));
    
    \ConfigStatusReg[17]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(17));
    
    \Stamp1ShadowReg2[15]\ : SLE
      port map(D => STAMP_0_data_frame(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(15));
    
    \APBState[0]\ : SLE
      port map(D => APBState_ns(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => APBState_Z(0));
    
    \StampFSMPC_6_0_a2[4]\ : CFG2
      generic map(INIT => x"2")

      port map(A => un8_tempcounter_cry_4_S, B => 
        ControllUnitState_Z(11), Y => StampFSMPC_6(4));
    
    \StampFSMR1[29]\ : SLE
      port map(D => pageaddr_5_i_m4(29), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(29));
    
    \readmemorylimitedcnt[0]\ : SLE
      port map(D => readmemorylimitedcnt_5(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorylimitedcnt_Z(0));
    
    \ReadMemoryState[2]\ : SLE
      port map(D => ReadMemoryState_Z(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ReadMemoryState_Z(2));
    
    \InternalData2Memory[31]\ : SLE
      port map(D => InternalData2Memory_27(31), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(31));
    
    \ControllUnitState[5]\ : SLE
      port map(D => ControllUnitState_ns(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(5));
    
    un1_currentaddrreg_cry_24 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(24), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_23_Z, S => 
        un1_currentaddrreg_cry_24_S, Y => 
        un1_currentaddrreg_cry_24_Y, FCO => 
        un1_currentaddrreg_cry_24_Z);
    
    \mainProcess.InternalData2Memory_27_0_iv_0[18]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(18), C => 
        Stamp1ShadowReg2_Z(18), D => 
        InternalData2Memory_27_0_iv_0_1(18), Y => 
        InternalData2Memory_27(18));
    
    \APB3ReadMemoryLimitedState_RNO[0]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => APB3ReadMemoryLimitedState_Z(2), B => 
        APB3ReadMemoryLimitedState_Z(4), C => N_50_0, D => 
        APB3ReadMemoryLimitedState_Z(3), Y => N_145_mux);
    
    \mainProcess.pageaddr_5_i_m4[8]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(8), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(8), Y => pageaddr_5_i_m4(8));
    
    \SPITransmitReg_RNO_1[14]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(14), Y => N_15_mux_16);
    
    \ControllUnitSubState_ns_i_a7_0[1]\ : CFG4
      generic map(INIT => x"A020")

      port map(A => ControllUnitSubState_ns_i_a7_0_2_Z(1), B => 
        ControllUnitState_Z(2), C => 
        ControllUnitSubState_ns_i_a7_0_3_Z(1), D => N_5700, Y => 
        N_2641);
    
    \ReadMemoryShadowReg[14]\ : SLE
      port map(D => InternalDataFromMem(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(14));
    
    \mainProcess.InternalAddr2Memory_34_m2[8]\ : CFG4
      generic map(INIT => x"AA8F")

      port map(A => InternalAddr2Memory_Z(8), B => 
        ControllUnitState_Z(11), C => 
        InternalAddr2Memory_34_m2_1_0(8), D => 
        InternalAddr2Memory_34_sm0, Y => 
        InternalAddr2Memory_34_m2(8));
    
    \un23_o3[1]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => ControllUnitState_Z(4), B => N_4343_i, C => 
        ControllUnitState_Z(7), Y => N_1262);
    
    \PRDATA[24]\ : SLE
      port map(D => PRDATA_8(24), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(24));
    
    \StampFSMR1[22]\ : SLE
      port map(D => pageaddr_5_i_m4(22), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(22));
    
    \StampFSMR1[11]\ : SLE
      port map(D => pageaddr_5_i_m4(11), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(11));
    
    \mainProcess.ConfigStatusReg_26_i_m2[31]\ : CFG4
      generic map(INIT => x"3AAA")

      port map(A => ConfigStatusReg_Z(31), B => SPIaddr_Z(0), C
         => ControllUnitState_Z(1), D => GPIO_6_M2F_c, Y => 
        N_4347);
    
    \mainProcess.PRDATA_8_0_iv_0[17]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(17), B => 
        PRDATA_8_0_iv_0_3(17), C => PRDATA_8_0_iv_0_6(17), Y => 
        PRDATA_8(17));
    
    \tempcounter[5]\ : SLE
      port map(D => N_4297_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_enabletimestampgen2_1_i, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tempcounter_Z(5));
    
    \SPITransmitReg[9]\ : SLE
      port map(D => SPITransmitReg_13(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(9));
    
    \Stamp1ShadowReg2[19]\ : SLE
      port map(D => STAMP_0_data_frame(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(19));
    
    \mainProcess.PRDATA_8_0_iv_0_1[10]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(2), B => CommandReg_Z(10), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(10));
    
    \mainProcess.PRDATA_8_0_iv_0_2[27]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(27), 
        D => CurrentAddrReg_Z(27), Y => PRDATA_8_0_iv_0_2(27));
    
    \ConfigStatusReg[30]\ : SLE
      port map(D => ConfigStatusReg_26(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ConfigStatusReg_Z(30));
    
    \APB3ReadMemoryLimitedState[5]\ : SLE
      port map(D => APB3ReadMemoryLimitedState_ns(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        APB3ReadMemoryLimitedState_Z(5));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[18]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(18), C => pageaddr(26), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(18));
    
    PRDATA_17_sqmuxa_2 : CFG4
      generic map(INIT => x"8000")

      port map(A => APBState_Z(0), B => sb_sb_0_STAMP_PADDR(3), C
         => sb_sb_0_STAMP_PADDR(2), D => sb_sb_0_STAMP_PADDR(6), 
        Y => PRDATA_17_sqmuxa_2_Z);
    
    \mainProcess.PRDATA_8_0_iv_0_1[3]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ConfigStatusReg_Z(3), B => CommandReg_Z(3), C
         => N_1025, D => N_4335, Y => PRDATA_8_0_iv_0_1(3));
    
    un8_tempcounter_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => StampFSMPC_Z(7), C => \GND\, D
         => \GND\, FCI => un8_tempcounter_cry_6_Z, S => 
        un8_tempcounter_cry_7_S, Y => un8_tempcounter_cry_7_Y, 
        FCO => un8_tempcounter_cry_7_Z);
    
    \SPITransmitReg_RNO_1[20]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(20), Y => N_15_mux_10);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[2]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(2), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(2));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[13]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(13), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0(13));
    
    \CommandReg[12]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(12));
    
    \mainProcess.SPITransmitReg_13_0_iv_0[3]\ : CFG4
      generic map(INIT => x"A808")

      port map(A => N_4270, B => InternalDataFromMem(3), C => 
        SPIState_1_sqmuxa, D => sb_sb_0_STAMP_PWDATA(3), Y => 
        SPITransmitReg_13(3));
    
    \ReadMemoryState_RNO[5]\ : CFG4
      generic map(INIT => x"0501")

      port map(A => N_80, B => ReadMemoryState_Z(5), C => 
        ReadMemoryState_ns_i_0_0_Z(3), D => N_2496, Y => N_2477_i);
    
    \Stamp1ShadowReg2[7]\ : SLE
      port map(D => STAMP_0_data_frame(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(7));
    
    \mainProcess.readmemorylimitedcnt_5[8]\ : CFG2
      generic map(INIT => x"2")

      port map(A => readmemorylimitedcnt_5_RNO_S(8), B => 
        APB3ReadMemoryLimitedState_Z(1), Y => 
        readmemorylimitedcnt_5(8));
    
    \InternalData2Memory[9]\ : SLE
      port map(D => InternalData2Memory_27(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(9));
    
    \InternalData2Memory[21]\ : SLE
      port map(D => InternalData2Memory_27(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(21));
    
    \ControllUnitState[2]\ : SLE
      port map(D => ControllUnitState_ns(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(2));
    
    \mainProcess.PRDATA_8_0_iv_0_1[12]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(4), B => CommandReg_Z(12), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(12));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[20]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(20), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(20));
    
    \SPITransmitReg_RNO_0[10]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(2), Y => N_4_21);
    
    \mainProcess.InternalAddr2Memory_34_14\ : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory_34_sm0, B => 
        InternalAddr2Memory_34_m0(3), C => N_143_mux, Y => 
        InternalAddr2Memory_34_14);
    
    \SPITransmitReg_RNO_1[17]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(17), Y => N_15_mux_13);
    
    \SPIState_RNIQS8J[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => SPIState_Z(3), B => SPIState_Z(1), Y => m46_0);
    
    \StampFSMR1[8]\ : SLE
      port map(D => pageaddr_5_i_m4(8), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(8));
    
    \mainProcess.PRDATA_8_0_iv_0_3[24]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(24), B => 
        Stamp1ShadowReg2_Z(24), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(24));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[19]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(19), C => pageaddr(27), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(19));
    
    \mainProcess.PRDATA_8_0_iv_0_1[13]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(5), B => CommandReg_Z(13), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(13));
    
    \APB3ReadMemoryLimitedState_RNIM0KJ[5]\ : CFG4
      generic map(INIT => x"0700")

      port map(A => APB3ReadMemoryLimitedState_Z(5), B => 
        ConfigStatusReg_Z(4), C => ControllUnitState_Z(13), D => 
        N_138, Y => N_143_mux);
    
    \readmemoryaddrcounter[30]\ : SLE
      port map(D => un1_readmemoryaddrcounter_cry_1_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \GND\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemoryaddrcounter_Z(30));
    
    \Stamp1ShadowReg1[8]\ : SLE
      port map(D => STAMP_0_data_frame(40), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(8));
    
    \readmemorylimitedcnt_RNI1LOJ[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemorylimitedcnt_Z(0), C => 
        \GND\, D => \GND\, FCI => 
        un1_readmemorylimitedcnt_cry_0_cy, S => 
        readmemorylimitedcnt_RNI1LOJ_S(0), Y => 
        readmemorylimitedcnt_RNI1LOJ_Y(0), FCO => 
        un1_readmemorylimitedcnt_cry_0);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[31]\ : CFG4
      generic map(INIT => x"ACA0")

      port map(A => SPIRecReg(31), B => pageaddr(7), C => 
        ReadMemoryState_Z(4), D => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(31));
    
    \Stamp1ShadowReg1[10]\ : SLE
      port map(D => STAMP_0_data_frame(42), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(10));
    
    \SPITransmitReg_RNO_1[8]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(8), Y => N_15_mux_22);
    
    \ConfigStatusReg_RNICDT61[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_2496_i, B => ConfigStatusReg_Z(4), Y => 
        N_81);
    
    \Stamp1ShadowReg1[31]\ : SLE
      port map(D => STAMP_0_data_frame(63), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(31));
    
    \mainProcess.InternalAddr2Memory_34_m0[2]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ControllUnitState_Z(2), B => 
        un1_memorycnt_1_cry_2_S, C => StampFSMPC_Z(2), Y => 
        InternalAddr2Memory_34_m0(2));
    
    \ReadMemoryShadowReg[26]\ : SLE
      port map(D => InternalDataFromMem(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(26));
    
    \SPITransmitReg_RNO[26]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_5, B => InternalDataFromMem(26), C => 
        N_54, D => N_15_mux_4, Y => SPITransmitReg_13(26));
    
    \ControllUnitState_RNI2VHT[14]\ : CFG3
      generic map(INIT => x"80")

      port map(A => ControllUnitState_Z(14), B => dataReady_0, C
         => GPIO_6_M2F_c, Y => ControllUnitState_RNI2VHT_Z(14));
    
    \SPITransmitReg_RNO[18]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_13, B => InternalDataFromMem(18), C => 
        N_54, D => N_15_mux_12, Y => SPITransmitReg_13(18));
    
    \CommandReg[6]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(6));
    
    GND_Z : GND
      port map(Y => \GND\);
    
    \mainProcess.PRDATA_8_0_iv_0_6[26]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(26), C => 
        PRDATA_8_0_iv_0_1(26), D => PRDATA_8_0_iv_0_0(26), Y => 
        PRDATA_8_0_iv_0_6(26));
    
    \mainProcess.PRDATA_8_0_iv_0_0[15]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(15), D => SPIRecReg(15), Y => 
        PRDATA_8_0_iv_0_0(15));
    
    \StampFSMR1[3]\ : SLE
      port map(D => pageaddr_5_i_m4(3), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(3));
    
    \ControllUnitSubState_ns_i_0[1]\ : CFG4
      generic map(INIT => x"4F0F")

      port map(A => InternalBusy, B => ControllUnitState_Z(2), C
         => N_4343, D => N_2648, Y => 
        ControllUnitSubState_ns_i_0_Z(1));
    
    un1_currentaddrreg_cry_22 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(22), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_21_Z, S => 
        un1_currentaddrreg_cry_22_S, Y => 
        un1_currentaddrreg_cry_22_Y, FCO => 
        un1_currentaddrreg_cry_22_Z);
    
    \SPITransmitReg[16]\ : SLE
      port map(D => SPITransmitReg_13(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(16));
    
    \ReadMemoryShadowReg[12]\ : SLE
      port map(D => InternalDataFromMem(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(12));
    
    \mainProcess.PRDATA_8_0_iv_0[8]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(8), B => 
        PRDATA_8_0_iv_0_3(8), C => PRDATA_8_0_iv_0_6(8), Y => 
        PRDATA_8(8));
    
    \mainProcess.pageaddr_5_i_m4[16]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(16), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(16), Y => pageaddr_5_i_m4(16));
    
    \SPITransmitReg_RNO_1[16]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(16), Y => N_15_mux_14);
    
    \mainProcess.PRDATA_8_0_iv_0_2[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(4), 
        D => CurrentAddrReg_Z(4), Y => PRDATA_8_0_iv_0_2(4));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[4]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(4), C => pageaddr(12), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(4));
    
    \ConfigStatusReg_RNO_1[3]\ : CFG4
      generic map(INIT => x"0104")

      port map(A => sb_sb_0_STAMP_PADDR(7), B => 
        ConfigStatusReg_Z(3), C => sb_sb_0_STAMP_PADDR(10), D => 
        sb_sb_0_STAMP_PWDATA(3), Y => m86_m7_0);
    
    \mainProcess.PRDATA_8_0_iv_0_3[19]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(19), B => 
        Stamp1ShadowReg2_Z(19), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(19));
    
    \un23_1[1]\ : CFG4
      generic map(INIT => x"FFE8")

      port map(A => ControllUnitState_Z(8), B => 
        ControllUnitSubState_Z(1), C => ControllUnitSubState_Z(0), 
        D => N_1298, Y => un23_1_Z(1));
    
    \ControllUnitState[12]\ : SLE
      port map(D => N_161, CLK => sb_sb_0_FIC_0_CLK, EN => 
        GPIO_6_M2F_c, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ControllUnitState_Z(12));
    
    \CurrentAddrReg[22]\ : SLE
      port map(D => un1_currentaddrreg_cry_22_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(22));
    
    \ControllUnitState_ns_0_0_a2_0[12]\ : CFG3
      generic map(INIT => x"20")

      port map(A => ControllUnitSubState_ns_i_a7_4_4_Z(1), B => 
        N_4339, C => ControllUnitSubState_ns_i_a7_4_5_Z(1), Y => 
        N_734);
    
    un1_memorycnt_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => memorycnt_Z(4), C => \GND\, D => 
        \GND\, FCI => un1_memorycnt_1_cry_3_Z, S => 
        un1_memorycnt_1_cry_4_S, Y => un1_memorycnt_1_cry_4_Y, 
        FCO => un1_memorycnt_1_cry_4_Z);
    
    StartAddrReg_0_sqmuxa_0_a2_0 : CFG4
      generic map(INIT => x"0080")

      port map(A => sb_sb_0_STAMP_PADDR(2), B => 
        sb_sb_0_STAMP_PADDR(5), C => sb_sb_0_STAMP_PADDR(4), D
         => sb_sb_0_STAMP_PADDR(3), Y => N_1029);
    
    \mainProcess.PRDATA_8_0_iv_0_0[5]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(5), D => SPIRecReg(5), Y => 
        PRDATA_8_0_iv_0_0(5));
    
    \tempcounter_RNO[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_1261_i, B => un8_tempcounter_cry_3_S, Y => 
        N_4295_i);
    
    \mainProcess.readmemorylimitedcnt_5[2]\ : CFG2
      generic map(INIT => x"2")

      port map(A => readmemorylimitedcnt_RNI4U3I1_S(2), B => 
        APB3ReadMemoryLimitedState_Z(1), Y => 
        readmemorylimitedcnt_5(2));
    
    \Command_RNIU9GL[4]\ : CFG2
      generic map(INIT => x"2")

      port map(A => Command_Z(0), B => Command_Z(4), Y => m33_e_0);
    
    \Stamp1ShadowReg1[22]\ : SLE
      port map(D => STAMP_0_data_frame(54), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(22));
    
    \SPITransmitReg_RNO_1[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_4272_i, B => ReadMemoryState_Z(8), Y => 
        SPITransmitReg_RNO_1_Z(0));
    
    \mainProcess.PRDATA_8_0_iv_0_6[15]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(15), C => 
        PRDATA_8_0_iv_0_1(15), D => PRDATA_8_0_iv_0_0(15), Y => 
        PRDATA_8_0_iv_0_6(15));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[12]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(12), B => 
        TimeStampValue(12), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(12));
    
    un1_readmemoryaddrcounter_cry_0 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemoryaddrcounter_Z(31), C
         => \GND\, D => \GND\, FCI => 
        un1_readmemoryaddrcounter_s_0_836_FCO, S => 
        un1_readmemoryaddrcounter_cry_0_S, Y => 
        un1_readmemoryaddrcounter_cry_0_Y, FCO => 
        un1_readmemoryaddrcounter_cry_0_Z);
    
    \SPITransmitReg[6]\ : SLE
      port map(D => SPITransmitReg_13(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(6));
    
    \mainProcess.InternalData2Memory_27_0_iv_1[13]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0(13), C => pageaddr(21), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_1(13));
    
    \InternalAddr2Memory[3]\ : SLE
      port map(D => InternalAddr2Memory_34(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => InternalAddr2Memory_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => InternalAddr2Memory_Z(3));
    
    \MemoryPageSize[7]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(7));
    
    \ReadMemoryShadowReg[1]\ : SLE
      port map(D => InternalDataFromMem(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(1));
    
    \StartAddrReg[17]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(17));
    
    \SPITransmitReg_RNO_0[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(1), Y => N_4_22);
    
    \PRDATA[20]\ : SLE
      port map(D => PRDATA_8(20), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(20));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[15]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(15), C => 
        Stamp1ShadowReg2_Z(15), D => 
        InternalData2Memory_27_0_iv_0_1(15), Y => 
        InternalData2Memory_27(15));
    
    \ControllUnitState_ns_i_0_a2_1_0[14]\ : CFG3
      generic map(INIT => x"01")

      port map(A => ControllUnitState_Z(2), B => 
        ControllUnitState_Z(0), C => ControllUnitState_Z(4), Y
         => ControllUnitState_ns_i_0_a2_1(14));
    
    \SPIState_RNO_1[2]\ : CFG4
      generic map(INIT => x"0C1D")

      port map(A => SPIState_Z(2), B => SPIState_Z(3), C => 
        N_150_mux, D => N_31_0, Y => SPIState_RNO_1_Z(2));
    
    \ReadMemoryShadowReg[18]\ : SLE
      port map(D => InternalDataFromMem(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(18));
    
    \mainProcess.InternalData2Memory_27_0_iv_1[25]\ : CFG4
      generic map(INIT => x"FCFA")

      port map(A => ControllUnitState_Z(11), B => SPIRecReg(25), 
        C => pageaddr_m(1), D => ReadMemoryState_Z(4), Y => 
        InternalData2Memory_27_0_iv_1(25));
    
    \mainProcess.InternalData2Memory_27_0_iv[13]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_3(13), C => 
        Stamp1ShadowReg2_Z(13), D => 
        InternalData2Memory_27_0_iv_1(13), Y => 
        InternalData2Memory_27(13));
    
    \mainProcess.PRDATA_8_0_iv_0_6[30]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(30), C => 
        PRDATA_8_0_iv_0_1(30), D => PRDATA_8_0_iv_0_0(30), Y => 
        PRDATA_8_0_iv_0_6(30));
    
    \StampFSMPC_6_0_a2[6]\ : CFG2
      generic map(INIT => x"2")

      port map(A => un8_tempcounter_cry_6_S, B => 
        ControllUnitState_Z(11), Y => StampFSMPC_6(6));
    
    SPIState_m2_e_1_1 : CFG4
      generic map(INIT => x"0004")

      port map(A => sb_sb_0_STAMP_PADDR(6), B => 
        sb_sb_0_STAMP_PADDR(5), C => sb_sb_0_STAMP_PADDR(8), D
         => sb_sb_0_STAMP_PADDR(9), Y => SPIState_m2_e_1_1_Z);
    
    InternalAddr2Memory_4_sqmuxa_i : CFG3
      generic map(INIT => x"7F")

      port map(A => ControllUnitState_Z(9), B => N_4343_i, C => 
        GPIO_6_M2F_c, Y => N_1232_i);
    
    \mainProcess.PRDATA_8_0_iv_0_1[14]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(6), B => CommandReg_Z(14), C
         => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(14));
    
    \mainProcess.InternalAddr2Memory_34_m0[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ControllUnitState_Z(2), B => 
        un1_memorycnt_1_cry_4_S, C => StampFSMPC_Z(4), Y => 
        InternalAddr2Memory_34_m0(4));
    
    \mainProcess.PRDATA_8_0_iv_0_3[4]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(4), B => 
        Stamp1ShadowReg2_Z(4), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(4));
    
    \StampFSMR1[21]\ : SLE
      port map(D => pageaddr_5_i_m4(21), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(21));
    
    \mainProcess.PRDATA_8_0_iv_0_0[27]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(27), D => SPIRecReg(27), Y => 
        PRDATA_8_0_iv_0_0(27));
    
    \InternalData2Memory[24]\ : SLE
      port map(D => InternalData2Memory_27(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(24));
    
    \ConfigStatusReg[22]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize(14));
    
    \SPITransmitReg[30]\ : SLE
      port map(D => SPITransmitReg_13(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(30));
    
    \APB3ReadMemoryLimitedState[3]\ : SLE
      port map(D => APB3ReadMemoryLimitedState_Z(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        APB3ReadMemoryLimitedState_Z(3));
    
    \tempcounter[4]\ : SLE
      port map(D => N_4296_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_enabletimestampgen2_1_i, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tempcounter_Z(4));
    
    \CurrentAddrReg[30]\ : SLE
      port map(D => un1_currentaddrreg_cry_30_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(30));
    
    \mainProcess.InternalAddr2Memory_34_m2s2\ : CFG2
      generic map(INIT => x"E")

      port map(A => ControllUnitState_Z(11), B => 
        ControllUnitState_Z(10), Y => InternalAddr2Memory_34_sm0);
    
    intRam : ram
      port map(InternalData2Memory(31) => 
        InternalData2Memory_Z(31), InternalData2Memory(30) => 
        InternalData2Memory_Z(30), InternalData2Memory(29) => 
        InternalData2Memory_Z(29), InternalData2Memory(28) => 
        InternalData2Memory_Z(28), InternalData2Memory(27) => 
        InternalData2Memory_Z(27), InternalData2Memory(26) => 
        InternalData2Memory_Z(26), InternalData2Memory(25) => 
        InternalData2Memory_Z(25), InternalData2Memory(24) => 
        InternalData2Memory_Z(24), InternalData2Memory(23) => 
        InternalData2Memory_Z(23), InternalData2Memory(22) => 
        InternalData2Memory_Z(22), InternalData2Memory(21) => 
        InternalData2Memory_Z(21), InternalData2Memory(20) => 
        InternalData2Memory_Z(20), InternalData2Memory(19) => 
        InternalData2Memory_Z(19), InternalData2Memory(18) => 
        InternalData2Memory_Z(18), InternalData2Memory(17) => 
        InternalData2Memory_Z(17), InternalData2Memory(16) => 
        InternalData2Memory_Z(16), InternalData2Memory(15) => 
        InternalData2Memory_Z(15), InternalData2Memory(14) => 
        InternalData2Memory_Z(14), InternalData2Memory(13) => 
        InternalData2Memory_Z(13), InternalData2Memory(12) => 
        InternalData2Memory_Z(12), InternalData2Memory(11) => 
        InternalData2Memory_Z(11), InternalData2Memory(10) => 
        InternalData2Memory_Z(10), InternalData2Memory(9) => 
        InternalData2Memory_Z(9), InternalData2Memory(8) => 
        InternalData2Memory_Z(8), InternalData2Memory(7) => 
        InternalData2Memory_Z(7), InternalData2Memory(6) => 
        InternalData2Memory_Z(6), InternalData2Memory(5) => 
        InternalData2Memory_Z(5), InternalData2Memory(4) => 
        InternalData2Memory_Z(4), InternalData2Memory(3) => 
        InternalData2Memory_Z(3), InternalData2Memory(2) => 
        InternalData2Memory_Z(2), InternalData2Memory(1) => 
        InternalData2Memory_Z(1), InternalData2Memory(0) => 
        InternalData2Memory_Z(0), InternalAddr2Memory(8) => 
        InternalAddr2Memory_Z(8), InternalAddr2Memory(7) => 
        InternalAddr2Memory_Z(7), InternalAddr2Memory(6) => 
        InternalAddr2Memory_Z(6), InternalAddr2Memory(5) => 
        InternalAddr2Memory_Z(5), InternalAddr2Memory(4) => 
        InternalAddr2Memory_Z(4), InternalAddr2Memory(3) => 
        InternalAddr2Memory_Z(3), InternalAddr2Memory(2) => 
        InternalAddr2Memory_Z(2), InternalAddr2Memory(1) => 
        InternalAddr2Memory_Z(1), InternalAddr2Memory(0) => 
        InternalAddr2Memory_Z(0), InternalDataFromMem(31) => 
        InternalDataFromMem(31), InternalDataFromMem(30) => 
        InternalDataFromMem(30), InternalDataFromMem(29) => 
        InternalDataFromMem(29), InternalDataFromMem(28) => 
        InternalDataFromMem(28), InternalDataFromMem(27) => 
        InternalDataFromMem(27), InternalDataFromMem(26) => 
        InternalDataFromMem(26), InternalDataFromMem(25) => 
        InternalDataFromMem(25), InternalDataFromMem(24) => 
        InternalDataFromMem(24), InternalDataFromMem(23) => 
        InternalDataFromMem(23), InternalDataFromMem(22) => 
        InternalDataFromMem(22), InternalDataFromMem(21) => 
        InternalDataFromMem(21), InternalDataFromMem(20) => 
        InternalDataFromMem(20), InternalDataFromMem(19) => 
        InternalDataFromMem(19), InternalDataFromMem(18) => 
        InternalDataFromMem(18), InternalDataFromMem(17) => 
        InternalDataFromMem(17), InternalDataFromMem(16) => 
        InternalDataFromMem(16), InternalDataFromMem(15) => 
        InternalDataFromMem(15), InternalDataFromMem(14) => 
        InternalDataFromMem(14), InternalDataFromMem(13) => 
        InternalDataFromMem(13), InternalDataFromMem(12) => 
        InternalDataFromMem(12), InternalDataFromMem(11) => 
        InternalDataFromMem(11), InternalDataFromMem(10) => 
        InternalDataFromMem(10), InternalDataFromMem(9) => 
        InternalDataFromMem(9), InternalDataFromMem(8) => 
        InternalDataFromMem(8), InternalDataFromMem(7) => 
        InternalDataFromMem(7), InternalDataFromMem(6) => 
        InternalDataFromMem(6), InternalDataFromMem(5) => 
        InternalDataFromMem(5), InternalDataFromMem(4) => 
        InternalDataFromMem(4), InternalDataFromMem(3) => 
        InternalDataFromMem(3), InternalDataFromMem(2) => 
        InternalDataFromMem(2), InternalDataFromMem(1) => 
        InternalDataFromMem(1), InternalDataFromMem(0) => 
        InternalDataFromMem(0), resetn => resetn, WriteEnable => 
        WriteEnable_Z, sb_sb_0_FIC_0_CLK => sb_sb_0_FIC_0_CLK, 
        resetn_arst => resetn_arst);
    
    SPITransmitReg_1_sqmuxa_2_i : CFG2
      generic map(INIT => x"B")

      port map(A => SPIState_1_sqmuxa, B => N_4270, Y => N_54);
    
    \Command_RNI9R801[7]\ : CFG3
      generic map(INIT => x"01")

      port map(A => Command_Z(7), B => Command_Z(6), C => 
        Command_Z(5), Y => m17_e_1);
    
    \mainProcess.pageaddr_5_i_m4[15]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(15), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(15), Y => pageaddr_5_i_m4(15));
    
    \PRDATA[23]\ : SLE
      port map(D => PRDATA_8(23), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(23));
    
    \SPITransmitReg_RNO[21]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_10, B => InternalDataFromMem(21), C => 
        N_54, D => N_15_mux_9, Y => SPITransmitReg_13(21));
    
    \StampFSMR1[18]\ : SLE
      port map(D => N_4370, CLK => sb_sb_0_FIC_0_CLK, EN => 
        ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        pageaddr(18));
    
    SPITransmitReg_0_sqmuxa_2_i_0 : CFG4
      generic map(INIT => x"ECFF")

      port map(A => GPIO_6_M2F_c, B => SPIState_1_sqmuxa, C => 
        un1_SPIState_8_0_a3_0_Z, D => N_4270, Y => N_16);
    
    \SPITransmitReg_RNO_0[21]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(13), Y => N_4_10);
    
    \Command[3]\ : SLE
      port map(D => N_174_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        Command_1_sqmuxa_1_i_Z, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        Command_Z(3));
    
    \ReadMemoryShadowReg[27]\ : SLE
      port map(D => InternalDataFromMem(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(27));
    
    \ReadMemoryState_ns_i_o4_RNIAVKO[0]\ : CFG3
      generic map(INIT => x"1D")

      port map(A => N_2496, B => SPIState_Z(4), C => Command_Z(0), 
        Y => m106_1_1);
    
    un1_currentaddrreg_cry_23 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(23), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_22_Z, S => 
        un1_currentaddrreg_cry_23_S, Y => 
        un1_currentaddrreg_cry_23_Y, FCO => 
        un1_currentaddrreg_cry_23_Z);
    
    \readmemorylimitedcnt_RNIF8HD1[1]\ : CFG3
      generic map(INIT => x"20")

      port map(A => readmemorylimitedcnt_Z(8), B => 
        readmemorylimitedcnt_Z(6), C => readmemorylimitedcnt_Z(1), 
        Y => m60_e_4);
    
    \APB3ReadMemoryLimitedState[1]\ : SLE
      port map(D => APB3ReadMemoryLimitedState_ns(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        APB3ReadMemoryLimitedState_Z(1));
    
    \mainProcess.memorycnt_6_cry_1_0\ : ARI1
      generic map(INIT => x"52122")

      port map(A => ControllUnitState_Z(3), B => memorycnt_Z(2), 
        C => ControllUnitState_RNI2VHT_Z(14), D => N_1255_i, FCI
         => memorycnt_6_cry_0, S => memorycnt_6(2), Y => 
        memorycnt_6_cry_1_0_Y, FCO => memorycnt_6_cry_1);
    
    \ControllUnitSubState_RNIDU3L[1]\ : CFG2
      generic map(INIT => x"B")

      port map(A => ControllUnitSubState_Z(0), B => 
        ControllUnitSubState_Z(1), Y => N_4339);
    
    \mainProcess.PRDATA_8_0_iv_0_6[28]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(28), C => 
        PRDATA_8_0_iv_0_1(28), D => PRDATA_8_0_iv_0_0(28), Y => 
        PRDATA_8_0_iv_0_6(28));
    
    un8_tempcounter_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => StampFSMPC_Z(6), C => \GND\, D
         => \GND\, FCI => un8_tempcounter_cry_5_Z, S => 
        un8_tempcounter_cry_6_S, Y => un8_tempcounter_cry_6_Y, 
        FCO => un8_tempcounter_cry_6_Z);
    
    un1_enabletimestampgen2_5_7 : CFG3
      generic map(INIT => x"FB")

      port map(A => un1_enabletimestampgen2_5_3_Z, B => N_1128, C
         => un1_enabletimestampgen2_5_2_Z, Y => 
        un1_enabletimestampgen2_5_7_Z);
    
    readmemorycounter_1_sqmuxa_1_i_o2 : CFG3
      generic map(INIT => x"FE")

      port map(A => ReadMemoryState_Z(8), B => 
        ReadMemoryState_Z(5), C => ReadMemoryState_Z(7), Y => 
        N_62);
    
    \mainProcess.InternalData2Memory_27_0_iv[29]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_2(29), C => 
        Stamp1ShadowReg2_Z(29), D => 
        InternalData2Memory_27_0_iv_0(29), Y => 
        InternalData2Memory_27(29));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[24]\ : CFG4
      generic map(INIT => x"ACA0")

      port map(A => SPIRecReg(24), B => pageaddr(0), C => 
        ReadMemoryState_Z(4), D => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0(24));
    
    \ConfigStatusReg[3]\ : SLE
      port map(D => N_87, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ConfigStatusReg_Z(3));
    
    \mainProcess.pageaddr_5_i_m4[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(6), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(6), Y => pageaddr_5_i_m4(6));
    
    \mainProcess.PRDATA_8_0_iv_0[23]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(23), B => 
        PRDATA_8_0_iv_0_3(23), C => PRDATA_8_0_iv_0_6(23), Y => 
        PRDATA_8(23));
    
    \mainProcess.memorycnt_6_cry_6\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => N_1541_i, C => N_2624_2, D => 
        \GND\, FCI => memorycnt_6_cry_5, S => memorycnt_6(7), Y
         => memorycnt_6_cry_6_Y, FCO => memorycnt_6_cry_6);
    
    \StartAddrReg[21]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(21));
    
    \ReadMemoryState_ns_i_m3_i[1]\ : CFG4
      generic map(INIT => x"CA0A")

      port map(A => ReadMemoryState_Z(8), B => 
        ReadMemoryState_Z(7), C => N_68, D => N_2496, Y => N_44);
    
    \mainProcess.InternalData2Memory_27_0_iv_0[31]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_2(31), C => 
        Stamp1ShadowReg2_Z(31), D => 
        InternalData2Memory_27_0_iv_0_0(31), Y => 
        InternalData2Memory_27(31));
    
    \mainProcess.PRDATA_8_0_iv_0_1[4]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ConfigStatusReg_Z(4), B => CommandReg_Z(4), C
         => N_1025, D => N_4335, Y => PRDATA_8_0_iv_0_1(4));
    
    \SPITransmitReg_RNO[17]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_14, B => InternalDataFromMem(17), C => 
        N_54, D => N_15_mux_13, Y => SPITransmitReg_13(17));
    
    \mainProcess.readmemorylimitedcnt_5[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => readmemorylimitedcnt_RNI29U21_S(1), B => 
        APB3ReadMemoryLimitedState_Z(1), Y => 
        readmemorylimitedcnt_5(1));
    
    \Stamp1ShadowReg2[10]\ : SLE
      port map(D => STAMP_0_data_frame(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(10));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[28]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(28), C => 
        Stamp1ShadowReg2_Z(28), D => 
        InternalData2Memory_27_0_iv_0_1(28), Y => 
        InternalData2Memory_27(28));
    
    \PRDATA[30]\ : SLE
      port map(D => PRDATA_8(30), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(30));
    
    \ControllUnitState_ns_i_0_a2_0_1_0[14]\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_765_1, B => N_1041, C => N_1185, Y => 
        ControllUnitState_ns_i_0_a2_0_1_Z(14));
    
    \CommandReg[3]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(3));
    
    \SPITransmitReg_RNO_1[24]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(24), Y => N_15_mux_6);
    
    \mainProcess.InternalAddr2Memory_34_m0[7]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ControllUnitState_Z(2), B => 
        un1_memorycnt_1_cry_7_S, C => StampFSMPC_Z(7), Y => 
        InternalAddr2Memory_34_m0(7));
    
    \mainProcess.PRDATA_8_0_iv_0_2[19]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(19), 
        D => CurrentAddrReg_Z(19), Y => PRDATA_8_0_iv_0_2(19));
    
    \ReadMemoryState_ns_i_o4_3_RNII5851[0]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => Command_Z(0), B => 
        ReadMemoryState_ns_i_o4_3_Z(0), C => Command_Z(6), D => 
        Command_Z(5), Y => N_2496_i);
    
    \PRDATA[11]\ : SLE
      port map(D => PRDATA_8(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(11));
    
    un1_currentaddrreg_cry_20 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(20), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_19_Z, S => 
        un1_currentaddrreg_cry_20_S, Y => 
        un1_currentaddrreg_cry_20_Y, FCO => 
        un1_currentaddrreg_cry_20_Z);
    
    \mainProcess.InternalAddr2Memory_34_m0[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ControllUnitState_Z(2), B => 
        un1_memorycnt_1_cry_3_S, C => StampFSMPC_Z(3), Y => 
        InternalAddr2Memory_34_m0(3));
    
    \Stamp1ShadowReg2[0]\ : SLE
      port map(D => STAMP_0_data_frame(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(0));
    
    \StampFSMR1[5]\ : SLE
      port map(D => pageaddr_5_i_m4(5), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(5));
    
    un1_readmemoryaddrcounter_s_0_836 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => ReadMemoryState_Z(4), C => \GND\, 
        D => \GND\, FCI => \VCC\, S => 
        un1_readmemoryaddrcounter_s_0_836_S, Y => 
        un1_readmemoryaddrcounter_s_0_836_Y, FCO => 
        un1_readmemoryaddrcounter_s_0_836_FCO);
    
    un1_currentaddrreg_cry_16 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => pageaddr(16), C => \GND\, D => 
        \GND\, FCI => un1_currentaddrreg_cry_15_Z, S => 
        un1_currentaddrreg_cry_16_S, Y => 
        un1_currentaddrreg_cry_16_Y, FCO => 
        un1_currentaddrreg_cry_16_Z);
    
    \ConfigStatusReg_RNO_0[29]\ : CFG4
      generic map(INIT => x"0FBB")

      port map(A => SPIState_ns(3), B => sb_sb_0_STAMP_PWDATA(29), 
        C => N_149_mux, D => N_4340, Y => m98_xx_mm_1);
    
    \mainProcess.readmemorylimitedcnt_5[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => readmemorylimitedcnt_RNI1LOJ_S(0), B => 
        APB3ReadMemoryLimitedState_Z(1), Y => 
        readmemorylimitedcnt_5(0));
    
    \CurrentAddrReg[10]\ : SLE
      port map(D => un1_currentaddrreg_cry_10_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(10));
    
    un1_SPIState_8_0_a3 : CFG2
      generic map(INIT => x"8")

      port map(A => enableSPI_0_sqmuxa_2, B => 
        un1_SPIState_8_0_a3_0_Z, Y => N_102);
    
    \ReadMemoryState_ns_i_0_a3_2_7[3]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => readmemoryaddrcounter_Z(31), B => 
        readmemoryaddrcounter_Z(29), C => 
        readmemoryaddrcounter_Z(28), D => 
        readmemoryaddrcounter_Z(26), Y => 
        ReadMemoryState_ns_i_0_a3_2_7_Z(3));
    
    \Stamp1ShadowReg1[25]\ : SLE
      port map(D => STAMP_0_data_frame(57), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(25));
    
    \SPIState_RNO_0[4]\ : CFG4
      generic map(INIT => x"FA8A")

      port map(A => m46_1_1_0_1, B => Command_Z(0), C => N_21_0, 
        D => m46_1_1_tz, Y => m46_1_1_0);
    
    \mainProcess.PRDATA_8_0_iv_0_6[0]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(0), C => 
        PRDATA_8_0_iv_0_1(0), D => PRDATA_8_0_iv_0_0(0), Y => 
        PRDATA_8_0_iv_0_6(0));
    
    \mainProcess.PRDATA_8_0_iv_0[12]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(12), B => 
        PRDATA_8_0_iv_0_3(12), C => PRDATA_8_0_iv_0_6(12), Y => 
        PRDATA_8(12));
    
    \mainProcess.pageaddr_5_i_m4[10]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(10), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(10), Y => pageaddr_5_i_m4(10));
    
    \SPITransmitReg_RNO_0[14]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(6), Y => N_4_17);
    
    \StartAddrReg[15]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(15));
    
    \StampFSMR1[10]\ : SLE
      port map(D => pageaddr_5_i_m4(10), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(10));
    
    \Stamp1ShadowReg1[3]\ : SLE
      port map(D => STAMP_0_data_frame(35), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(3));
    
    \mainProcess.PRDATA_8_0_iv_0_0[10]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(10), D => SPIRecReg(10), Y => 
        PRDATA_8_0_iv_0_0(10));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[23]\ : CFG4
      generic map(INIT => x"FEEE")

      port map(A => N_4527, B => 
        InternalData2Memory_27_0_iv_0_1(23), C => SPIRecReg(23), 
        D => ReadMemoryState_Z(4), Y => 
        InternalData2Memory_27(23));
    
    \mainProcess.InternalData2Memory_27_0_iv_2[26]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(26), B => 
        TimeStampValue(26), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_2(26));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[6]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(6), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(6));
    
    \mainProcess.pageaddr_5_i_m4[14]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(14), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(14), Y => pageaddr_5_i_m4(14));
    
    \readmemorycounter_RNO_0[3]\ : CFG4
      generic map(INIT => x"0B0F")

      port map(A => N_4268, B => un1_enableSPI_1_sqmuxa_1_i, C
         => readmemorycounter_Z(3), D => readmemorycounter_Z(2), 
        Y => N_95);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[4]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(4), B => TimeStampValue(4), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(4));
    
    un1_currentaddrreg_cry_14 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize(14), B => pageaddr(14), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_13_Z, S
         => un1_currentaddrreg_cry_14_S, Y => 
        un1_currentaddrreg_cry_14_Y, FCO => 
        un1_currentaddrreg_cry_14_Z);
    
    \ConfigStatusReg[31]\ : SLE
      port map(D => N_249_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => ConfigStatusReg_Z(31));
    
    \mainProcess.InternalData2Memory_27_0_iv_2[27]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(27), B => 
        TimeStampValue(27), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_2(27));
    
    \mainProcess.InternalAddr2Memory_34[8]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => InternalAddr2Memory_34_m2(8), B => 
        InternalAddr2Memory_34_m5(8), C => N_143_mux, Y => 
        InternalAddr2Memory_34(8));
    
    \InternalData2Memory[22]\ : SLE
      port map(D => InternalData2Memory_27(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(22));
    
    \ControllUnitState[14]\ : SLE
      port map(D => ControllUnitState_ns(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \GND\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(14));
    
    \CommandReg[1]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(1));
    
    \SPITransmitReg_RNO[12]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_19, B => InternalDataFromMem(12), C => 
        N_54, D => N_15_mux_18, Y => SPITransmitReg_13(12));
    
    \mainProcess.PRDATA_8_0_iv_0[21]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(21), B => 
        PRDATA_8_0_iv_0_3(21), C => PRDATA_8_0_iv_0_6(21), Y => 
        PRDATA_8(21));
    
    \mainProcess.InternalAddr2Memory_34_m2_1_1[0]\ : CFG3
      generic map(INIT => x"5C")

      port map(A => StampFSMPC_Z(0), B => 
        ControllUnitSubState_Z(0), C => ControllUnitState_Z(2), Y
         => InternalAddr2Memory_34_m2_1_1(0));
    
    \Command[4]\ : SLE
      port map(D => N_172_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        Command_1_sqmuxa_1_i_Z, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        Command_Z(4));
    
    InternalData2Memory_0_sqmuxa_1_i : CFG2
      generic map(INIT => x"7")

      port map(A => N_4343_i, B => ControllUnitState_Z(8), Y => 
        N_1128);
    
    \ControllUnitState[0]\ : SLE
      port map(D => N_2554_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        GPIO_6_M2F_c, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ControllUnitState_Z(0));
    
    \Stamp1ShadowReg2[22]\ : SLE
      port map(D => STAMP_0_data_frame(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(22));
    
    \Stamp1ShadowReg1[29]\ : SLE
      port map(D => STAMP_0_data_frame(61), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(29));
    
    \SPITransmitReg_RNO_1[31]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(31), Y => N_15_mux);
    
    \ReadMemoryState_ns_i_o4[0]\ : CFG4
      generic map(INIT => x"FFFD")

      port map(A => Command_Z(0), B => 
        ReadMemoryState_ns_i_o4_3_Z(0), C => Command_Z(6), D => 
        Command_Z(5), Y => N_2496);
    
    \readmemorylimitedcnt_RNI7K912[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemorylimitedcnt_Z(3), C => 
        \GND\, D => \GND\, FCI => un1_readmemorylimitedcnt_cry_2, 
        S => readmemorylimitedcnt_RNI7K912_S(3), Y => 
        readmemorylimitedcnt_RNI7K912_Y(3), FCO => 
        un1_readmemorylimitedcnt_cry_3);
    
    \SPITransmitReg_RNO_1[27]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(27), Y => N_15_mux_3);
    
    \mainProcess.PRDATA_8_0_iv_0_1[0]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ConfigStatusReg_Z(0), B => CommandReg_Z(0), C
         => N_1025, D => N_4335, Y => PRDATA_8_0_iv_0_1(0));
    
    \mainProcess.memorycnt_6_cry_5\ : ARI1
      generic map(INIT => x"48800")

      port map(A => \VCC\, B => N_1541_i, C => memorycnt_Z(6), D
         => \GND\, FCI => memorycnt_6_cry_4, S => memorycnt_6(6), 
        Y => memorycnt_6_cry_5_Y, FCO => memorycnt_6_cry_5);
    
    \Stamp1ShadowReg2[30]\ : SLE
      port map(D => STAMP_0_data_frame(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(30));
    
    un1_currentaddrreg_cry_7 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(7), B => pageaddr(7), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_6_Z, S
         => un1_currentaddrreg_cry_7_S, Y => 
        un1_currentaddrreg_cry_7_Y, FCO => 
        un1_currentaddrreg_cry_7_Z);
    
    \SPIState[4]\ : SLE
      port map(D => N_157_mux, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => SPIState_Z(4));
    
    \mainProcess.PRDATA_8_0_iv_0_0[1]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(1), D => SPIRecReg(1), Y => 
        PRDATA_8_0_iv_0_0(1));
    
    \mainProcess.PRDATA_8_0_iv_0_0[12]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(12), D => SPIRecReg(12), Y => 
        PRDATA_8_0_iv_0_0(12));
    
    \tempcounter_RNO[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_1261_i, B => un8_tempcounter_cry_2_S, Y => 
        N_139_i);
    
    \mainProcess.PRDATA_8_0_iv_0_2[25]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(25), 
        D => CurrentAddrReg_Z(25), Y => PRDATA_8_0_iv_0_2(25));
    
    \InternalData2Memory[4]\ : SLE
      port map(D => InternalData2Memory_27(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(4));
    
    \mainProcess.PRDATA_8_0_iv_0_6[10]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(10), C => 
        PRDATA_8_0_iv_0_1(10), D => PRDATA_8_0_iv_0_0(10), Y => 
        PRDATA_8_0_iv_0_6(10));
    
    \InternalData2Memory[10]\ : SLE
      port map(D => InternalData2Memory_27(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(10));
    
    \ControllUnitState_ns_i_0_a4[14]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => ControllUnitState_Z(2), B => N_765_1, C => 
        N_4339, D => N_4349, Y => N_765);
    
    \mainProcess.PRDATA_8_0_iv_0[25]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(25), B => 
        PRDATA_8_0_iv_0_3(25), C => PRDATA_8_0_iv_0_6(25), Y => 
        PRDATA_8(25));
    
    \SPITransmitReg[5]\ : SLE
      port map(D => SPITransmitReg_13(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(5));
    
    \Stamp1ShadowReg2[8]\ : SLE
      port map(D => STAMP_0_data_frame(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(8));
    
    \mainProcess.PRDATA_8_0_iv_0_3[5]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(5), B => 
        Stamp1ShadowReg2_Z(5), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(5));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[0]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(0), C => 
        Stamp1ShadowReg2_Z(0), D => 
        InternalData2Memory_27_0_iv_0_1(0), Y => 
        InternalData2Memory_27(0));
    
    \SPITransmitReg[19]\ : SLE
      port map(D => SPITransmitReg_13(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(19));
    
    \StartAddrReg[29]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(29));
    
    \mainProcess.PRDATA_8_0_iv_0_0[13]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(13), D => SPIRecReg(13), Y => 
        PRDATA_8_0_iv_0_0(13));
    
    \mainProcess.pageaddr_5_i_m4[0]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(0), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(0), Y => pageaddr_5_i_m4(0));
    
    \SPITransmitReg[23]\ : SLE
      port map(D => SPITransmitReg_13(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(23));
    
    \mainProcess.readmemorycounter_6_iv[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => N_4259, B => N_4254_i, Y => 
        readmemorycounter_6(1));
    
    \SPITransmitReg_RNO_0[17]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(9), Y => N_4_14);
    
    \mainProcess.InternalData2Memory_27_0_iv_1_RNO[25]\ : CFG3
      generic map(INIT => x"40")

      port map(A => ReadMemoryState_Z(4), B => pageaddr(1), C => 
        ControllUnitState_Z(10), Y => pageaddr_m(1));
    
    \ReadMemoryState_ns_0_a3_0_a3[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_68, B => ReadMemoryState_Z(5), Y => 
        ReadMemoryState_ns(4));
    
    un1_SPIState_8_0_a3_0 : CFG2
      generic map(INIT => x"2")

      port map(A => enableSPI_1_sqmuxa_1_0_Z, B => InternalBusy, 
        Y => un1_SPIState_8_0_a3_0_Z);
    
    \SPITransmitReg_RNO[0]\ : CFG4
      generic map(INIT => x"FBFA")

      port map(A => N_13_mux_1, B => N_54, C => 
        SPITransmitReg_RNO_1_Z(0), D => InternalDataFromMem(0), Y
         => SPITransmitReg_13(0));
    
    \APB3ReadMemoryLimitedState_RNO[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_139_mux, B => 
        APB3ReadMemoryLimitedState_Z(3), Y => 
        APB3ReadMemoryLimitedState_ns(4));
    
    \mainProcess.InternalAddr2Memory_34_m0[5]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ControllUnitState_Z(2), B => 
        un1_memorycnt_1_cry_5_S, C => StampFSMPC_Z(5), Y => 
        InternalAddr2Memory_34_m0(5));
    
    \ControllUnitState_ns_i_a2[11]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => memorycnt_Z(4), B => memorycnt_Z(8), C => 
        N_2624_1, D => ControllUnitState_ns_i_a2_3_Z(11), Y => 
        N_2624);
    
    \ControllUnitState[8]\ : SLE
      port map(D => ControllUnitState_ns(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(8));
    
    \mainProcess.PRDATA_8_0_iv_0_6[21]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(21), C => 
        PRDATA_8_0_iv_0_1(21), D => PRDATA_8_0_iv_0_0(21), Y => 
        PRDATA_8_0_iv_0_6(21));
    
    \mainProcess.PRDATA_8_0_iv_0_6[12]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(12), C => 
        PRDATA_8_0_iv_0_1(12), D => PRDATA_8_0_iv_0_0(12), Y => 
        PRDATA_8_0_iv_0_6(12));
    
    \readmemorylimitedcnt_RNI4U3I1[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemorylimitedcnt_Z(2), C => 
        \GND\, D => \GND\, FCI => un1_readmemorylimitedcnt_cry_1, 
        S => readmemorylimitedcnt_RNI4U3I1_S(2), Y => 
        readmemorylimitedcnt_RNI4U3I1_Y(2), FCO => 
        un1_readmemorylimitedcnt_cry_2);
    
    \PRDATA[25]\ : SLE
      port map(D => PRDATA_8(25), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(25));
    
    \ControllUnitState[13]\ : SLE
      port map(D => N_7_0, CLK => sb_sb_0_FIC_0_CLK, EN => 
        GPIO_6_M2F_c, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ControllUnitState_Z(13));
    
    \ReadMemoryShadowReg[29]\ : SLE
      port map(D => InternalDataFromMem(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(29));
    
    \mainProcess.pageaddr_5[27]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(27), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(27), Y => pageaddr_5(27));
    
    \ControllUnitState_RNO[13]\ : CFG2
      generic map(INIT => x"8")

      port map(A => dataReady_0, B => ControllUnitState_Z(14), Y
         => N_7_0);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[8]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(8), C => pageaddr(16), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(8));
    
    \memorycnt[1]\ : SLE
      port map(D => memorycnt_6_cry_0_0_Y, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \GND\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        memorycnt_Z(1));
    
    \mainProcess.PRDATA_8_0_iv_0[3]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => PRDATA_8_0_iv_0_2(3), B => 
        PRDATA_8_0_iv_0_3(3), C => PRDATA_8_0_iv_0_6(3), Y => 
        PRDATA_8(3));
    
    \mainProcess.InternalAddr2Memory_34[5]\ : CFG4
      generic map(INIT => x"FDDD")

      port map(A => InternalAddr2Memory_34_1(5), B => 
        InternalAddr2Memory_34_2, C => 
        readmemoryaddrcounter_Z(26), D => ReadMemoryState_Z(4), Y
         => InternalAddr2Memory_34(5));
    
    \mainProcess.PRDATA_8_0_iv_0_6[13]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(13), C => 
        PRDATA_8_0_iv_0_1(13), D => PRDATA_8_0_iv_0_0(13), Y => 
        PRDATA_8_0_iv_0_6(13));
    
    \Stamp1ShadowReg1[17]\ : SLE
      port map(D => STAMP_0_data_frame(49), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(17));
    
    \StartAddrReg[28]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(28));
    
    \CommandReg[25]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(25));
    
    \mainProcess.PRDATA_8_0_iv_0_3[2]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(2), B => 
        Stamp1ShadowReg2_Z(2), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(2));
    
    \SPITransmitReg_RNO_1[26]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(26), Y => N_15_mux_4);
    
    \mainProcess.PRDATA_8_0_iv_0_3[16]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(16), B => 
        Stamp1ShadowReg2_Z(16), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(16));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[22]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(22), B => 
        TimeStampValue(22), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(22));
    
    \mainProcess.PRDATA_8_0_iv_0_2[1]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(1), 
        D => CurrentAddrReg_Z(1), Y => PRDATA_8_0_iv_0_2(1));
    
    \un23_o3_i_o4[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => ControllUnitSubState_Z(0), B => 
        ControllUnitSubState_Z(1), Y => N_4343);
    
    \mainProcess.pageaddr_5_i_m4[22]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(22), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(22), Y => pageaddr_5_i_m4(22));
    
    \ConfigStatusReg_RNO[3]\ : CFG4
      generic map(INIT => x"55B4")

      port map(A => ReadMemoryState_Z(3), B => 
        ConfigStatusReg_Z(3), C => m86_0_1, D => N_2496_i, Y => 
        N_87);
    
    \SPITransmitReg_RNO[8]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_23, B => InternalDataFromMem(8), C => 
        N_54, D => N_15_mux_22, Y => SPITransmitReg_13(8));
    
    \ConfigStatusReg[5]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(5));
    
    \Stamp1ShadowReg2[4]\ : SLE
      port map(D => STAMP_0_data_frame(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(4));
    
    \SPITransmitReg_RNO[24]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => N_4_7, B => InternalDataFromMem(24), C => 
        N_54, D => N_15_mux_6, Y => SPITransmitReg_13(24));
    
    \mainProcess.InternalAddr2Memory_34_1[4]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => readmemorylimitedcnt_Z(4), B => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), C => N_138, Y
         => InternalAddr2Memory_34_1(4));
    
    \CurrentAddrReg[14]\ : SLE
      port map(D => un1_currentaddrreg_cry_14_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(14));
    
    \StartAddrReg[7]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(7));
    
    \Stamp1ShadowReg1[13]\ : SLE
      port map(D => STAMP_0_data_frame(45), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(13));
    
    \PRDATA[0]\ : SLE
      port map(D => PRDATA_8(0), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(0));
    
    \mainProcess.PRDATA_8_0_iv_0_3[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(29), B => 
        Stamp1ShadowReg2_Z(29), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(29));
    
    \readmemoryaddrcounter_3[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => ReadMemoryState_ns(5), B => 
        un1_readmemoryaddrcounter_s_8_S, Y => 
        readmemoryaddrcounter_3_Z(8));
    
    \StampFSMR1[28]\ : SLE
      port map(D => pageaddr_5_i_m4(28), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(28));
    
    \ControllUnitState_RNO[3]\ : CFG4
      generic map(INIT => x"0F0D")

      port map(A => N_2624, B => ControllUnitState_Z(4), C => 
        ControllUnitState_ns_i_0_2_Z(11), D => N_4339, Y => 
        N_2550_i);
    
    \ControllUnitState_ns_0_0_o2[12]\ : CFG2
      generic map(INIT => x"D")

      port map(A => ControllUnitSubState_Z(0), B => 
        ControllUnitSubState_Z(1), Y => N_4342);
    
    \ControllUnitState[4]\ : SLE
      port map(D => ControllUnitState_ns(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => GPIO_6_M2F_c, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ControllUnitState_Z(4));
    
    \SPITransmitReg_RNO_0[16]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(8), Y => N_4_15);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[16]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(16), B => 
        TimeStampValue(16), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(16));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[7]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(7), C => pageaddr(15), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(7));
    
    \SPITransmitReg_RNO_1[11]\ : CFG3
      generic map(INIT => x"80")

      port map(A => SPIState_1_sqmuxa, B => N_4270, C => 
        sb_sb_0_STAMP_PWDATA(11), Y => N_15_mux_19);
    
    \MemoryPageSize[11]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(11));
    
    un1_currentaddrreg_cry_12 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(12), B => pageaddr(12), C
         => \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_11_Z, 
        S => un1_currentaddrreg_cry_12_S, Y => 
        un1_currentaddrreg_cry_12_Y, FCO => 
        un1_currentaddrreg_cry_12_Z);
    
    un1_currentaddrreg_cry_4 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(4), B => pageaddr(4), C => 
        \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_3_Z, S
         => un1_currentaddrreg_cry_4_S, Y => 
        un1_currentaddrreg_cry_4_Y, FCO => 
        un1_currentaddrreg_cry_4_Z);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[2]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(2), C => pageaddr(10), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(2));
    
    \readmemorylimitedcnt_RNI29U21[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemorylimitedcnt_Z(1), C => 
        \GND\, D => \GND\, FCI => un1_readmemorylimitedcnt_cry_0, 
        S => readmemorylimitedcnt_RNI29U21_S(1), Y => 
        readmemorylimitedcnt_RNI29U21_Y(1), FCO => 
        un1_readmemorylimitedcnt_cry_1);
    
    un1_readmemoryaddrcounter_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => readmemoryaddrcounter_Z(24), C
         => \GND\, D => \GND\, FCI => 
        un1_readmemoryaddrcounter_cry_6_Z, S => 
        un1_readmemoryaddrcounter_cry_7_S, Y => 
        un1_readmemoryaddrcounter_cry_7_Y, FCO => 
        un1_readmemoryaddrcounter_cry_7_Z);
    
    \ConfigStatusReg_RNIM7LI[0]\ : CFG4
      generic map(INIT => x"6000")

      port map(A => ConfigStatusReg_Z(0), B => 
        ConfigStatusReg_Z(1), C => GPIO_6_M2F_c, D => 
        ControllUnitState_Z(13), Y => N_4294_i);
    
    \Command_RNI4K1M2[4]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => Command_Z(0), B => N_21_0, C => Command_Z(4), 
        Y => N_71);
    
    \mainProcess.PRDATA_8_0_iv_0_1[27]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ConfigStatusReg_Z(27), B => CommandReg_Z(27), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(27));
    
    \ControllUnitSubState_ns_0_0_a2_1[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => ControllUnitState_Z(1), B => 
        ControllUnitState_Z(10), C => ControllUnitState_Z(12), D
         => ControllUnitState_Z(0), Y => N_1035);
    
    \Stamp1ShadowReg2[25]\ : SLE
      port map(D => STAMP_0_data_frame(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(25));
    
    \ReadMemoryState[5]\ : SLE
      port map(D => N_2477_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => ReadMemoryState_Z(5));
    
    \mainProcess.readmemorylimitedcnt_5[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => readmemorylimitedcnt_RNIG3LV2_S(5), B => 
        APB3ReadMemoryLimitedState_Z(1), Y => 
        readmemorylimitedcnt_5(5));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[4]\ : CFG4
      generic map(INIT => x"FFEC")

      port map(A => InternalData2Memory_5_sqmuxa_Z, B => 
        InternalData2Memory_27_0_iv_0_3(4), C => 
        Stamp1ShadowReg2_Z(4), D => 
        InternalData2Memory_27_0_iv_0_1(4), Y => 
        InternalData2Memory_27(4));
    
    \CommandReg[15]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => Command_1_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => CommandReg_Z(15));
    
    \Stamp1ShadowReg2[9]\ : SLE
      port map(D => STAMP_0_data_frame(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(9));
    
    \ConfigStatusReg[2]\ : SLE
      port map(D => N_88, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ConfigStatusReg_Z(2));
    
    \Stamp1ShadowReg2[6]\ : SLE
      port map(D => STAMP_0_data_frame(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(6));
    
    TimeStampGen : Timestamp
      port map(TimeStampValue(31) => TimeStampValue(31), 
        TimeStampValue(30) => TimeStampValue(30), 
        TimeStampValue(29) => TimeStampValue(29), 
        TimeStampValue(28) => TimeStampValue(28), 
        TimeStampValue(27) => TimeStampValue(27), 
        TimeStampValue(26) => TimeStampValue(26), 
        TimeStampValue(25) => TimeStampValue(25), 
        TimeStampValue(24) => TimeStampValue(24), 
        TimeStampValue(23) => TimeStampValue(23), 
        TimeStampValue(22) => TimeStampValue(22), 
        TimeStampValue(21) => TimeStampValue(21), 
        TimeStampValue(20) => TimeStampValue(20), 
        TimeStampValue(19) => TimeStampValue(19), 
        TimeStampValue(18) => TimeStampValue(18), 
        TimeStampValue(17) => TimeStampValue(17), 
        TimeStampValue(16) => TimeStampValue(16), 
        TimeStampValue(15) => TimeStampValue(15), 
        TimeStampValue(14) => TimeStampValue(14), 
        TimeStampValue(13) => TimeStampValue(13), 
        TimeStampValue(12) => TimeStampValue(12), 
        TimeStampValue(11) => TimeStampValue(11), 
        TimeStampValue(10) => TimeStampValue(10), 
        TimeStampValue(9) => TimeStampValue(9), TimeStampValue(8)
         => TimeStampValue(8), TimeStampValue(7) => 
        TimeStampValue(7), TimeStampValue(6) => TimeStampValue(6), 
        TimeStampValue(5) => TimeStampValue(5), TimeStampValue(4)
         => TimeStampValue(4), TimeStampValue(3) => 
        TimeStampValue(3), TimeStampValue(2) => TimeStampValue(2), 
        TimeStampValue(1) => TimeStampValue(1), TimeStampValue(0)
         => TimeStampValue(0), getTime => getTime_Z, 
        enableTimestampGen => enableTimestampGen_Z, 
        sb_sb_0_FIC_0_CLK => sb_sb_0_FIC_0_CLK, resetn_arst => 
        resetn_arst);
    
    Command_1_sqmuxa_1_i : CFG3
      generic map(INIT => x"F8")

      port map(A => m73_m2_e_2, B => Command_1_sqmuxa_0_a2_0_Z, C
         => SPIState_RNI27U44_Z(1), Y => Command_1_sqmuxa_1_i_Z);
    
    \mainProcess.InternalAddr2Memory_34_m5[8]\ : CFG4
      generic map(INIT => x"C0A0")

      port map(A => readmemoryaddrcounter_Z(23), B => 
        readmemorylimitedcnt_Z(8), C => N_4266, D => N_138, Y => 
        InternalAddr2Memory_34_m5(8));
    
    PRDATA_17_sqmuxa : CFG4
      generic map(INIT => x"0200")

      port map(A => PRDATA_17_sqmuxa_8_Z, B => 
        un1_APBState_1_2_0_Z, C => sb_sb_0_STAMP_PADDR(11), D => 
        PRDATA_17_sqmuxa_2_Z, Y => PRDATA_17_sqmuxa_Z);
    
    \Stamp1ShadowReg1[16]\ : SLE
      port map(D => STAMP_0_data_frame(48), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(16));
    
    \ControllUnitState_ns_i_0_a2_3[14]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => ControllUnitState_Z(6), B => N_4351, C => 
        ControllUnitState_Z(8), D => ControllUnitState_Z(9), Y
         => N_1185);
    
    \PRDATA[9]\ : SLE
      port map(D => PRDATA_8(9), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(9));
    
    un1_APBState_1_1 : CFG3
      generic map(INIT => x"FB")

      port map(A => \un1_APBState_1_5_1z\, B => APBState_Z(0), C
         => sb_sb_0_STAMP_PADDR(11), Y => un1_APBState_1_1_Z);
    
    un1_currentaddrreg_cry_0 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize(0), B => pageaddr(0), C => 
        \GND\, D => \GND\, FCI => \GND\, S => 
        un1_currentaddrreg_cry_0_S, Y => 
        un1_currentaddrreg_cry_0_Y, FCO => 
        un1_currentaddrreg_cry_0_Z);
    
    \PRDATA[8]\ : SLE
      port map(D => PRDATA_8(8), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(8));
    
    \mainProcess.PRDATA_8_0_iv_0_0[14]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(14), D => SPIRecReg(14), Y => 
        PRDATA_8_0_iv_0_0(14));
    
    \ControllUnitState_RNI8UAF[12]\ : CFG2
      generic map(INIT => x"8")

      port map(A => GPIO_6_M2F_c, B => ControllUnitState_Z(12), Y
         => N_1080_i);
    
    \mainProcess.InternalAddr2Memory_34_m4_i[0]\ : CFG2
      generic map(INIT => x"7")

      port map(A => ReadMemoryState_Z(4), B => 
        readmemoryaddrcounter_Z(31), Y => N_4258);
    
    \Stamp1ShadowReg2[29]\ : SLE
      port map(D => STAMP_0_data_frame(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(29));
    
    \CurrentAddrReg[16]\ : SLE
      port map(D => un1_currentaddrreg_cry_16_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(16));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_1[6]\ : CFG4
      generic map(INIT => x"DCCC")

      port map(A => ReadMemoryState_Z(4), B => 
        InternalData2Memory_27_0_iv_0_0(6), C => pageaddr(14), D
         => ControllUnitState_Z(11), Y => 
        InternalData2Memory_27_0_iv_0_1(6));
    
    \InternalData2Memory[13]\ : SLE
      port map(D => InternalData2Memory_27(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(13));
    
    \StampFSMR1[20]\ : SLE
      port map(D => pageaddr_5_i_m4(20), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(20));
    
    \mainProcess.ConfigStatusReg_26_0_1[30]\ : CFG4
      generic map(INIT => x"0DFF")

      port map(A => ControllUnitSubState_Z(1), B => N_2624, C => 
        N_4343_i, D => ConfigStatusReg_26_0_a2_1(30), Y => 
        ConfigStatusReg_26_0_1(30));
    
    \CurrentAddrReg[0]\ : SLE
      port map(D => un1_currentaddrreg_cry_0_Y, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(0));
    
    \mainProcess.InternalData2Memory_27_0_iv_2[29]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(29), B => 
        TimeStampValue(29), C => InternalData2Memory_4_sqmuxa_Z, 
        D => InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_2(29));
    
    \mainProcess.ConfigStatusReg_26_0[30]\ : CFG4
      generic map(INIT => x"3FAA")

      port map(A => sb_sb_0_STAMP_PWDATA(30), B => 
        ConfigStatusReg_26_0_m2_1(30), C => 
        ConfigStatusReg_26_0_1(30), D => N_4340, Y => 
        ConfigStatusReg_26(30));
    
    \ControllUnitState_ns_i_0_0[14]\ : CFG4
      generic map(INIT => x"B333")

      port map(A => ControllUnitState_ns_i_0_a2_1(14), B => 
        ConfigStatusReg_Z(2), C => N_1185, D => N_4350, Y => 
        ControllUnitState_ns_i_0_0_Z(14));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(0), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(0));
    
    InternalAddr2Memory_4_sqmuxa_i_o3 : CFG2
      generic map(INIT => x"7")

      port map(A => N_4343_i, B => ControllUnitState_Z(9), Y => 
        N_1254);
    
    \StampFSMR1[9]\ : SLE
      port map(D => pageaddr_5_i_m4(9), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(9));
    
    \Stamp1ShadowReg2[3]\ : SLE
      port map(D => STAMP_0_data_frame(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(3));
    
    \PRDATA[22]\ : SLE
      port map(D => PRDATA_8(22), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(22));
    
    \ControllUnitState_ns_0_0_a2_1[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_4339, B => ConfigStatusReg_Z(2), Y => 
        N_1045);
    
    \ControllUnitState_ns_0_0[10]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => ControllUnitState_Z(5), B => 
        ControllUnitState_Z(4), C => N_4339, D => N_1045, Y => 
        ControllUnitState_ns(10));
    
    \ControllUnitState_ns_0[6]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ControllUnitState_Z(9), B => 
        ControllUnitState_Z(8), C => N_1045, D => N_4339, Y => 
        ControllUnitState_ns(6));
    
    \mainProcess.PRDATA_8_0_iv_0_2[20]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(20), 
        D => CurrentAddrReg_Z(20), Y => PRDATA_8_0_iv_0_2(20));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_3[9]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => Stamp1ShadowReg1_Z(9), B => TimeStampValue(9), 
        C => InternalData2Memory_4_sqmuxa_Z, D => 
        InternalData2Memory_3_sqmuxa_Z, Y => 
        InternalData2Memory_27_0_iv_0_3(9));
    
    \mainProcess.InternalAddr2Memory_34_10\ : CFG3
      generic map(INIT => x"40")

      port map(A => InternalAddr2Memory_34_sm0, B => 
        InternalAddr2Memory_34_m0(7), C => N_143_mux, Y => 
        InternalAddr2Memory_34_10);
    
    \mainProcess.ConfigStatusReg_26_0_o2[30]\ : CFG4
      generic map(INIT => x"2FFF")

      port map(A => N_1316_i, B => ControllUnitState_Z(14), C => 
        GPIO_6_M2F_c, D => ConfigStatusReg_24_sn_N_5, Y => N_4354);
    
    \mainProcess.PRDATA_8_0_iv_0_0[31]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(31), D => SPIRecReg(31), Y => 
        PRDATA_8_0_iv_0_0(31));
    
    \PRDATA[29]\ : SLE
      port map(D => PRDATA_8(29), CLK => sb_sb_0_FIC_0_CLK, EN
         => un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(29));
    
    \mainProcess.PRDATA_8_0_iv_0_6[14]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => N_1033, B => Stamp1ShadowReg1_Z(14), C => 
        PRDATA_8_0_iv_0_1(14), D => PRDATA_8_0_iv_0_0(14), Y => 
        PRDATA_8_0_iv_0_6(14));
    
    \CurrentAddrReg[9]\ : SLE
      port map(D => un1_currentaddrreg_cry_9_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(9));
    
    \mainProcess.PRDATA_8_0_iv_0_0[25]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => un1_paddr_3, B => N_1031, C => 
        ReadMemoryShadowReg_Z(25), D => SPIRecReg(25), Y => 
        PRDATA_8_0_iv_0_0(25));
    
    \un23_i_a2_0[0]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => ControllUnitState_Z(5), B => 
        ControllUnitState_Z(6), C => ControllUnitSubState_Z(1), D
         => N_1041, Y => N_762);
    
    \Stamp1ShadowReg1[1]\ : SLE
      port map(D => STAMP_0_data_frame(33), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(1));
    
    \InternalData2Memory[15]\ : SLE
      port map(D => InternalData2Memory_27(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(15));
    
    \CurrentAddrReg[31]\ : SLE
      port map(D => un1_currentaddrreg_cry_30_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(31));
    
    \CurrentAddrReg[28]\ : SLE
      port map(D => un1_currentaddrreg_cry_28_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(28));
    
    \mainProcess.PRDATA_8_0_iv_0_3[18]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(18), B => 
        Stamp1ShadowReg2_Z(18), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(18));
    
    \InternalData2Memory[29]\ : SLE
      port map(D => InternalData2Memory_27(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(29));
    
    \InternalData2Memory[26]\ : SLE
      port map(D => InternalData2Memory_27(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(26));
    
    \mainProcess.PRDATA_8_0_iv_0_2[8]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(8), 
        D => CurrentAddrReg_Z(8), Y => PRDATA_8_0_iv_0_2(8));
    
    InternalAddr2Memory_0_sqmuxa_0 : CFG2
      generic map(INIT => x"1")

      port map(A => ReadMemoryState_Z(4), B => 
        ReadMemoryState_Z(3), Y => N_138);
    
    \MemoryPageSize[4]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => MemoryPageSize_Z(4));
    
    \tempcounter_RNO[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_1261_i, B => un8_tempcounter_cry_4_S, Y => 
        N_4296_i);
    
    \CurrentAddrReg[23]\ : SLE
      port map(D => un1_currentaddrreg_cry_23_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(23));
    
    \ReadMemoryShadowReg[15]\ : SLE
      port map(D => InternalDataFromMem(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => ReadMemoryShadowReg_0_sqmuxa_i_Z, 
        ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => ReadMemoryShadowReg_Z(15));
    
    \mainProcess.PRDATA_8_0_iv_0_2[16]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(16), 
        D => CurrentAddrReg_Z(16), Y => PRDATA_8_0_iv_0_2(16));
    
    \mainProcess.pageaddr_5_i_m4[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(2), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(2), Y => pageaddr_5_i_m4(2));
    
    \ControllUnitSubState_ns_i_a7_4_3[1]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => memorycnt_Z(8), B => memorycnt_Z(4), C => 
        memorycnt_Z(3), D => N_2624_2, Y => 
        ControllUnitSubState_ns_i_a7_4_3_Z(1));
    
    \ConfigStatusReg_RNO_2[29]\ : CFG4
      generic map(INIT => x"0454")

      port map(A => ControllUnitState_Z(1), B => N_89, C => N_146, 
        D => SPIState_ns(3), Y => m94_1_1);
    
    un1_currentaddrreg_cry_13 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(13), B => pageaddr(13), C
         => \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_12_Z, 
        S => un1_currentaddrreg_cry_13_S, Y => 
        un1_currentaddrreg_cry_13_Y, FCO => 
        un1_currentaddrreg_cry_13_Z);
    
    \tempcounter_RNO[6]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_1261_i, B => un8_tempcounter_cry_6_S, Y => 
        N_4298_i);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[3]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(3), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(3));
    
    \mainProcess.PRDATA_8_0_iv_0_2[22]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(22), 
        D => CurrentAddrReg_Z(22), Y => PRDATA_8_0_iv_0_2(22));
    
    \mainProcess.pageaddr_5_i_m4[21]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => CurrentAddrReg_Z(21), B => isfirstrun_Z(0), C
         => StartAddrReg_Z(21), Y => pageaddr_5_i_m4(21));
    
    \ConfigStatusReg[26]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4340_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => ConfigStatusReg_Z(26));
    
    \mainProcess.InternalAddr2Memory_34[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => InternalAddr2Memory_34_m5(1), B => 
        InternalAddr2Memory_34_m2(1), C => N_143_mux, Y => 
        InternalAddr2Memory_34(1));
    
    \ConfigStatusReg[1]\ : SLE
      port map(D => N_252_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => resetn_arst, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => ConfigStatusReg_Z(1));
    
    \SPIState_RNO_5[2]\ : CFG3
      generic map(INIT => x"19")

      port map(A => N_21_0, B => SPIState_Z(4), C => Command_Z(0), 
        Y => SPIState_RNO_5_Z(2));
    
    un1_ControllUnitState_9_0 : CFG2
      generic map(INIT => x"D")

      port map(A => N_1254, B => ControllUnitState_Z(11), Y => 
        un1_ControllUnitState_9);
    
    \APB3ReadMemoryLimitedState_RNO[5]\ : CFG3
      generic map(INIT => x"E0")

      port map(A => APB3ReadMemoryLimitedState_Z(0), B => 
        APB3ReadMemoryLimitedState_Z(2), C => PRDATA_17_sqmuxa_Z, 
        Y => APB3ReadMemoryLimitedState_ns(0));
    
    PRDATA_17_sqmuxa_8 : CFG4
      generic map(INIT => x"0001")

      port map(A => sb_sb_0_STAMP_PADDR(0), B => 
        sb_sb_0_STAMP_PADDR(1), C => sb_sb_0_STAMP_PADDR(5), D
         => sb_sb_0_STAMP_PADDR(4), Y => PRDATA_17_sqmuxa_8_Z);
    
    \mainProcess.PRDATA_8_0_iv_0_1[19]\ : CFG4
      generic map(INIT => x"CE0A")

      port map(A => MemoryPageSize_Z(11), B => CommandReg_Z(19), 
        C => N_4335, D => N_1025, Y => PRDATA_8_0_iv_0_1(19));
    
    \SPITransmitReg_RNO_0[25]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1034, B => CommandReg_Z(17), Y => N_4_6);
    
    \SPITransmitReg[28]\ : SLE
      port map(D => SPITransmitReg_13(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_16, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        SPITransmitReg_Z(28));
    
    \mainProcess.PRDATA_8_0_iv_0_2[23]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_1032, B => N_1029, C => StartAddrReg_Z(23), 
        D => CurrentAddrReg_Z(23), Y => PRDATA_8_0_iv_0_2(23));
    
    un1_enableSPI_1_sqmuxa_1_0_0 : CFG4
      generic map(INIT => x"CE0A")

      port map(A => N_62, B => ReadMemoryState_Z(6), C => 
        N_4272_i, D => N_4274, Y => un1_enableSPI_1_sqmuxa_1_i);
    
    \Stamp1ShadowReg2[17]\ : SLE
      port map(D => STAMP_0_data_frame(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(17));
    
    \SPIState_RNO_4[2]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => Command_Z(0), B => SPIState_Z(4), C => 
        N_2496_i, D => N_21_0, Y => N_31_0);
    
    \Stamp1ShadowReg1[20]\ : SLE
      port map(D => STAMP_0_data_frame(52), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg1_Z(20));
    
    \StartAddrReg[2]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(2));
    
    \mainProcess.InternalData2Memory_27_0_iv_0[30]\ : CFG4
      generic map(INIT => x"ACA0")

      port map(A => SPIRecReg(30), B => pageaddr(6), C => 
        ReadMemoryState_Z(4), D => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0(30));
    
    enableSPI : SLE
      port map(D => un1_SPIState_8, CLK => sb_sb_0_FIC_0_CLK, EN
         => enableSPI_0_sqmuxa_3_i_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        enable);
    
    \tempcounter_RNO[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_1261_i, B => un8_tempcounter_s_8_S, Y => 
        N_4299_i);
    
    \readmemorylimitedcnt[3]\ : SLE
      port map(D => readmemorylimitedcnt_5(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorylimitedcnt_Z(3));
    
    \mainProcess.SPITransmitReg_13_0_iv_0[7]\ : CFG4
      generic map(INIT => x"A808")

      port map(A => N_4270, B => InternalDataFromMem(7), C => 
        SPIState_1_sqmuxa, D => sb_sb_0_STAMP_PWDATA(7), Y => 
        SPITransmitReg_13(7));
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[12]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(12), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(12));
    
    \InternalData2Memory[5]\ : SLE
      port map(D => InternalData2Memory_27(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        InternalData2Memory_0_sqmuxa_6_i_Z, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => InternalData2Memory_Z(5));
    
    \mainProcess.PRDATA_8_0_iv_0_1[30]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => ConfigStatusReg_Z(30), B => CommandReg_Z(30), 
        C => N_1025, D => N_4335, Y => PRDATA_8_0_iv_0_1(30));
    
    un1_currentaddrreg_cry_10 : ARI1
      generic map(INIT => x"555AA")

      port map(A => MemoryPageSize_Z(10), B => pageaddr(10), C
         => \GND\, D => \GND\, FCI => un1_currentaddrreg_cry_9_Z, 
        S => un1_currentaddrreg_cry_10_S, Y => 
        un1_currentaddrreg_cry_10_Y, FCO => 
        un1_currentaddrreg_cry_10_Z);
    
    \ControllUnitSubState_ns_i_a7_4_5[1]\ : CFG3
      generic map(INIT => x"20")

      port map(A => ControllUnitState_Z(3), B => 
        ControllUnitSubState_Z(0), C => 
        ControllUnitSubState_ns_i_a7_4_3_Z(1), Y => 
        ControllUnitSubState_ns_i_a7_4_5_Z(1));
    
    \mainProcess.getTime_3_f0\ : CFG4
      generic map(INIT => x"CCC4")

      port map(A => N_1254, B => N_1128, C => getTime_Z, D => 
        ControllUnitState_Z(10), Y => getTime_3);
    
    \StampFSMPC_6_0_a2[7]\ : CFG2
      generic map(INIT => x"2")

      port map(A => un8_tempcounter_cry_7_S, B => 
        ControllUnitState_Z(11), Y => StampFSMPC_6(7));
    
    \mainProcess.tempcounter_7_iv_i[7]\ : CFG3
      generic map(INIT => x"32")

      port map(A => N_1261_i, B => ControllUnitState_Z(1), C => 
        un8_tempcounter_cry_7_S, Y => tempcounter_7_iv_i(7));
    
    \StartAddrReg[8]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => StartAddrReg_0_sqmuxa, ALn => 
        resetn_arst, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => StartAddrReg_Z(8));
    
    \mainProcess.InternalAddr2Memory_34_ss3_i_0_m2\ : CFG3
      generic map(INIT => x"CA")

      port map(A => ReadMemoryState_Z(4), B => 
        APB3ReadMemoryLimitedState_RNI12J4_Y(5), C => N_138, Y
         => N_4266);
    
    \Stamp1ShadowReg2[13]\ : SLE
      port map(D => STAMP_0_data_frame(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_1080_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => Stamp1ShadowReg2_Z(13));
    
    \ControllUnitSubState_ns_i_a7_0_3[1]\ : CFG3
      generic map(INIT => x"10")

      port map(A => ControllUnitState_Z(5), B => 
        ControllUnitState_Z(6), C => N_1041, Y => 
        ControllUnitSubState_ns_i_a7_0_3_Z(1));
    
    \isfirstrun[0]\ : SLE
      port map(D => \VCC\, CLK => sb_sb_0_FIC_0_CLK, EN => 
        isfirstrun_1_sqmuxa, ALn => resetn_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        isfirstrun_Z(0));
    
    \mainProcess.PRDATA_8_0_iv_0_3[3]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => SPITransmitReg_Z(3), B => 
        Stamp1ShadowReg2_Z(3), C => N_1030, D => N_1026, Y => 
        PRDATA_8_0_iv_0_3(3));
    
    un1_ReadMemoryState_12_0_a2_0_a3 : CFG2
      generic map(INIT => x"1")

      port map(A => N_62, B => ReadMemoryState_Z(6), Y => 
        N_1508_i);
    
    \CurrentAddrReg[11]\ : SLE
      port map(D => un1_currentaddrreg_cry_11_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_4294_i, ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => CurrentAddrReg_Z(11));
    
    \StampFSMR1[14]\ : SLE
      port map(D => pageaddr_5_i_m4(14), CLK => sb_sb_0_FIC_0_CLK, 
        EN => ControllUnitState_RNI2VHT_Z(14), ALn => resetn_arst, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => pageaddr(14));
    
    \readmemorylimitedcnt[7]\ : SLE
      port map(D => readmemorylimitedcnt_5(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => resetn_arst, ADn
         => \GND\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        readmemorylimitedcnt_Z(7));
    
    \PRDATA[4]\ : SLE
      port map(D => PRDATA_8(4), CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_APBState_1_i, ALn => resetn_arst, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_Memory_PRDATA(4));
    
    MemoryPageSize_1_sqmuxa_0_o4 : CFG4
      generic map(INIT => x"FFFD")

      port map(A => PRDATA_17_sqmuxa_8_Z, B => 
        un1_APBState_1_2_0_Z, C => sb_sb_0_STAMP_PADDR(11), D => 
        MemoryPageSize_1_sqmuxa_0_o4_0_Z, Y => N_4340);
    
    \APB3ReadMemoryLimitedState_RNO[2]\ : CFG4
      generic map(INIT => x"0C2E")

      port map(A => APB3ReadMemoryLimitedState_Z(2), B => 
        APB3ReadMemoryLimitedState_Z(3), C => N_139_mux, D => 
        PRDATA_17_sqmuxa_Z, Y => N_101);
    
    WriteEnable : SLE
      port map(D => N_4265_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        WriteEnable_0_sqmuxa_i_Z, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        WriteEnable_Z);
    
    \mainProcess.InternalData2Memory_27_0_iv_0_0[4]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => ReadMemoryState_Z(4), B => SPIRecReg(4), C
         => ControllUnitState_Z(10), Y => 
        InternalData2Memory_27_0_iv_0_0(4));
    
    \ControllUnitState[3]\ : SLE
      port map(D => N_2550_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        GPIO_6_M2F_c, ALn => resetn_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => 
        ControllUnitState_Z(3));
    
    \tempcounter[2]\ : SLE
      port map(D => N_139_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_enabletimestampgen2_1_i, ALn => resetn_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        tempcounter_Z(2));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sb_sb_MSS is

    port( sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : in    std_logic_vector(31 downto 0);
          dataReady_0                             : in    std_logic;
          sb_sb_0_STAMP_PWDATA                    : out   std_logic_vector(31 downto 0);
          STAMP_PADDRS                            : out   std_logic_vector(15 downto 12);
          sb_sb_0_STAMP_PADDR                     : out   std_logic_vector(11 downto 0);
          sb_sb_0_FIC_0_CLK                       : in    std_logic;
          RXSM_SODS_c                             : in    std_logic;
          RXSM_SOE_c                              : in    std_logic;
          RXSM_LO_c                               : in    std_logic;
          FIC_0_LOCK                              : in    std_logic;
          PREADY_N_7                              : in    std_logic;
          PRDATA_N_5_i                            : in    std_logic;
          GPIO_6_M2F_c                            : out   std_logic;
          LED_RECORDING_c                         : out   std_logic;
          LED_HEARTBEAT_c                         : out   std_logic;
          sb_sb_0_STAMP_PWRITE                    : out   std_logic;
          sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx  : out   std_logic;
          sb_sb_0_STAMP_PENABLE                   : out   std_logic;
          sb_sb_0_GPIO_4_M2F                      : out   std_logic;
          sb_sb_0_GPIO_3_M2F                      : out   std_logic;
          DAPI_RX                                 : in    std_logic;
          DAPI_TX                                 : out   std_logic;
          TM_RX                                   : in    std_logic;
          TM_TX                                   : out   std_logic
        );

end sb_sb_MSS;

architecture DEF_ARCH of sb_sb_MSS is 

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component MSS_010

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component TRIBUFF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal EDAC_ERROR : std_logic_vector(7 downto 0);
    signal F_FM0_RDATA : std_logic_vector(31 downto 0);
    signal FIC_0_APB_M_PADDR : std_logic_vector(31 downto 16);
    signal F_HM0_SIZE : std_logic_vector(1 downto 0);
    signal FAB_OPMODE : std_logic_vector(1 downto 0);
    signal FAB_VCONTROL : std_logic_vector(3 downto 0);
    signal FAB_XCVRSEL : std_logic_vector(1 downto 0);
    signal FAB_XDATAOUT : std_logic_vector(7 downto 0);
    signal FIC32_0_MASTER : std_logic_vector(1 downto 0);
    signal FIC32_1_MASTER : std_logic_vector(1 downto 0);
    signal H2F_INTERRUPT : std_logic_vector(15 downto 0);
    signal FIC_2_APB_M_PADDR : std_logic_vector(15 downto 2);
    signal FIC_2_APB_M_PWDATA : std_logic_vector(31 downto 0);
    signal TCGF : std_logic_vector(9 downto 0);
    signal TRACEDATA : std_logic_vector(3 downto 0);
    signal TXD_RIF : std_logic_vector(3 downto 0);
    signal TXDF : std_logic_vector(7 downto 0);
    signal F_BID : std_logic_vector(3 downto 0);
    signal F_BRESP_HRESP0 : std_logic_vector(1 downto 0);
    signal F_RDATA_HRDATA01 : std_logic_vector(63 downto 0);
    signal F_RID : std_logic_vector(3 downto 0);
    signal F_RRESP_HRESP1 : std_logic_vector(1 downto 0);
    signal MDDR_FABRIC_PRDATA : std_logic_vector(15 downto 0);
    signal DRAM_ADDR : std_logic_vector(15 downto 0);
    signal DRAM_BA : std_logic_vector(2 downto 0);
    signal DRAM_DM_RDQS_OUT : std_logic_vector(2 downto 0);
    signal DRAM_DQ_OUT : std_logic_vector(17 downto 0);
    signal DRAM_DQS_OUT : std_logic_vector(2 downto 0);
    signal DRAM_FIFO_WE_OUT : std_logic_vector(1 downto 0);
    signal DM_OE : std_logic_vector(2 downto 0);
    signal DRAM_DQ_OE : std_logic_vector(17 downto 0);
    signal DRAM_DQS_OE : std_logic_vector(2 downto 0);
    signal MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        MMUART_1_RXD_PAD_Y, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, 
        MMUART_0_RXD_PAD_Y, CAN_RXBUS_MGPIO3A_H2F_A, 
        CAN_TX_EBL_MGPIO4A_H2F_A, CAN_TXBUS_MGPIO2A_H2F_A, 
        CAN_TXBUS_MGPIO2A_H2F_B, FIC_2_APB_M_PCLK, COMMS_INT, 
        FIC_2_APB_M_PRESET_N, F_FM0_READYOUT, F_FM0_RESP, 
        F_HM0_TRANS1, FAB_CHRGVBUS, FAB_DISCHRGVBUS, 
        FAB_DMPULLDOWN, FAB_DPPULLDOWN, FAB_DRVVBUS, FAB_IDPULLUP, 
        FAB_SUSPENDM, FAB_TERMSEL, FAB_TXVALID, FAB_VCONTROLLOADM, 
        FACC_GLMUX_SEL, MSS_RESET_N_M2F, GTX_CLK, H2F_NMI, 
        H2FCALIB, I2C0_SCL_MGPIO31B_H2F_A, 
        I2C0_SDA_MGPIO30B_H2F_A, I2C1_SCL_MGPIO1A_H2F_A, 
        I2C1_SCL_MGPIO1A_H2F_B, I2C1_SDA_MGPIO0A_H2F_A, 
        I2C1_SDA_MGPIO0A_H2F_B, MDCF, MDOENF, MDOF, 
        MMUART0_CTS_MGPIO19B_H2F_A, MMUART0_CTS_MGPIO19B_H2F_B, 
        MMUART0_DCD_MGPIO22B_H2F_A, MMUART0_DCD_MGPIO22B_H2F_B, 
        MMUART0_DSR_MGPIO20B_H2F_A, MMUART0_DSR_MGPIO20B_H2F_B, 
        MMUART0_DTR_MGPIO18B_H2F_A, MMUART0_DTR_MGPIO18B_H2F_B, 
        MMUART0_RI_MGPIO21B_H2F_A, MMUART0_RI_MGPIO21B_H2F_B, 
        MMUART0_RTS_MGPIO17B_H2F_A, MMUART0_RTS_MGPIO17B_H2F_B, 
        MMUART0_RXD_MGPIO28B_H2F_A, MMUART0_RXD_MGPIO28B_H2F_B, 
        MMUART0_SCK_MGPIO29B_H2F_A, MMUART0_SCK_MGPIO29B_H2F_B, 
        MMUART0_TXD_MGPIO27B_H2F_A, MMUART0_TXD_MGPIO27B_H2F_B, 
        MMUART1_DTR_MGPIO12B_H2F_A, MMUART1_RTS_MGPIO11B_H2F_A, 
        MMUART1_RTS_MGPIO11B_H2F_B, MMUART1_RXD_MGPIO26B_H2F_A, 
        MMUART1_RXD_MGPIO26B_H2F_B, MMUART1_SCK_MGPIO25B_H2F_A, 
        MMUART1_SCK_MGPIO25B_H2F_B, MMUART1_TXD_MGPIO24B_H2F_A, 
        MMUART1_TXD_MGPIO24B_H2F_B, MPLL_LOCK, 
        FIC_2_APB_M_PENABLE, FIC_2_APB_M_PSEL, FIC_2_APB_M_PWRITE, 
        RTC_MATCH, SLEEPDEEP, SLEEPHOLDACK, SLEEPING, 
        SMBALERT_NO0, SMBALERT_NO1, SMBSUS_NO0, SMBSUS_NO1, 
        SPI0_CLK_OUT, SPI0_SDI_MGPIO5A_H2F_A, 
        SPI0_SDI_MGPIO5A_H2F_B, SPI0_SDO_MGPIO6A_H2F_A, 
        SPI0_SS0_MGPIO7A_H2F_A, SPI0_SS0_MGPIO7A_H2F_B, 
        SPI0_SS1_MGPIO8A_H2F_A, SPI0_SS1_MGPIO8A_H2F_B, 
        SPI0_SS2_MGPIO9A_H2F_A, SPI0_SS2_MGPIO9A_H2F_B, 
        SPI0_SS3_MGPIO10A_H2F_A, SPI0_SS3_MGPIO10A_H2F_B, 
        SPI0_SS4_MGPIO19A_H2F_A, SPI0_SS5_MGPIO20A_H2F_A, 
        SPI0_SS6_MGPIO21A_H2F_A, SPI0_SS7_MGPIO22A_H2F_A, 
        SPI1_CLK_OUT, SPI1_SDI_MGPIO11A_H2F_A, 
        SPI1_SDI_MGPIO11A_H2F_B, SPI1_SDO_MGPIO12A_H2F_A, 
        SPI1_SDO_MGPIO12A_H2F_B, SPI1_SS0_MGPIO13A_H2F_A, 
        SPI1_SS0_MGPIO13A_H2F_B, SPI1_SS1_MGPIO14A_H2F_A, 
        SPI1_SS1_MGPIO14A_H2F_B, SPI1_SS2_MGPIO15A_H2F_A, 
        SPI1_SS2_MGPIO15A_H2F_B, SPI1_SS3_MGPIO16A_H2F_A, 
        SPI1_SS3_MGPIO16A_H2F_B, SPI1_SS4_MGPIO17A_H2F_A, 
        SPI1_SS5_MGPIO18A_H2F_A, SPI1_SS6_MGPIO23A_H2F_A, 
        SPI1_SS7_MGPIO24A_H2F_A, TRACECLK, TX_CLK, TX_ENF, 
        TX_ERRF, TXCTL_EN_RIF, TXEV, WDOGTIMEOUT, 
        F_ARREADY_HREADYOUT1, F_AWREADY_HREADYOUT0, F_BVALID, 
        F_RLAST, F_RVALID, F_WREADY, MDDR_FABRIC_PREADY, 
        MDDR_FABRIC_PSLVERR, \VCC\, \GND\, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT, DRAM_CASN, DRAM_CKE, 
        DRAM_CLK, DRAM_CSN, DRAM_ODT, DRAM_RASN, DRAM_RSTN, 
        DRAM_WEN, I2C0_SCL_USBC_DATA1_MGPIO31B_OUT, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OUT, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT, 
        MMUART0_DCD_MGPIO22B_OUT, MMUART0_DSR_MGPIO20B_OUT, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT, 
        MMUART0_RI_MGPIO21B_OUT, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT, 
        RGMII_MDC_RMII_MDC_OUT, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT, RGMII_RX_CLK_OUT, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT, 
        RGMII_RXD3_USBB_DATA4_OUT, RGMII_TX_CLK_OUT, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT, 
        RGMII_TXD2_USBB_DATA5_OUT, RGMII_TXD3_USBB_DATA6_OUT, 
        SPI0_SCK_USBA_XCLK_OUT, SPI0_SDI_USBA_DIR_MGPIO5A_OUT, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT, SPI1_SCK_OUT, 
        SPI1_SDI_MGPIO11A_OUT, SPI1_SDO_MGPIO12A_OUT, 
        SPI1_SS0_MGPIO13A_OUT, SPI1_SS1_MGPIO14A_OUT, 
        SPI1_SS2_MGPIO15A_OUT, SPI1_SS3_MGPIO16A_OUT, 
        SPI1_SS4_MGPIO17A_OUT, SPI1_SS5_MGPIO18A_OUT, 
        SPI1_SS6_MGPIO23A_OUT, SPI1_SS7_MGPIO24A_OUT, 
        USBC_XCLK_OUT, CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE, 
        MMUART0_DCD_MGPIO22B_OE, MMUART0_DSR_MGPIO20B_OE, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OE, 
        MMUART0_RI_MGPIO21B_OE, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE, 
        RGMII_MDC_RMII_MDC_OE, RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE, 
        RGMII_RX_CLK_OE, RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE, 
        RGMII_RXD3_USBB_DATA4_OE, RGMII_TX_CLK_OE, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE, 
        RGMII_TXD2_USBB_DATA5_OE, RGMII_TXD3_USBB_DATA6_OE, 
        SPI0_SCK_USBA_XCLK_OE, SPI0_SDI_USBA_DIR_MGPIO5A_OE, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE, SPI1_SCK_OE, 
        SPI1_SDI_MGPIO11A_OE, SPI1_SDO_MGPIO12A_OE, 
        SPI1_SS0_MGPIO13A_OE, SPI1_SS1_MGPIO14A_OE, 
        SPI1_SS2_MGPIO15A_OE, SPI1_SS3_MGPIO16A_OE, 
        SPI1_SS4_MGPIO17A_OE, SPI1_SS5_MGPIO18A_OE, 
        SPI1_SS6_MGPIO23A_OE, SPI1_SS7_MGPIO24A_OE, USBC_XCLK_OE
         : std_logic;

begin 


    MMUART_0_RXD_PAD : INBUF
      generic map(IOSTD => "")

      port map(PAD => DAPI_RX, Y => MMUART_0_RXD_PAD_Y);
    
    MSS_ADLIB_INST : MSS_010

              generic map(INIT => "00" & x"0000000003612000000000000000036100080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFF82FAF09007C33C804000006092C0000003FFFFE4000000000020100000000F0F01C000001825F84010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem",
         RTC_MAIN_XTL_FREQ => 0.000000, RTC_MAIN_XTL_MODE => "",
         DDR_CLK_FREQ => 100.000000)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => CAN_RXBUS_MGPIO3A_H2F_A, 
        CAN_RXBUS_MGPIO3A_H2F_B => sb_sb_0_GPIO_3_M2F, 
        CAN_TX_EBL_MGPIO4A_H2F_A => CAN_TX_EBL_MGPIO4A_H2F_A, 
        CAN_TX_EBL_MGPIO4A_H2F_B => sb_sb_0_GPIO_4_M2F, 
        CAN_TXBUS_MGPIO2A_H2F_A => CAN_TXBUS_MGPIO2A_H2F_A, 
        CAN_TXBUS_MGPIO2A_H2F_B => CAN_TXBUS_MGPIO2A_H2F_B, 
        CLK_CONFIG_APB => FIC_2_APB_M_PCLK, COMMS_INT => 
        COMMS_INT, CONFIG_PRESET_N => FIC_2_APB_M_PRESET_N, 
        EDAC_ERROR(7) => EDAC_ERROR(7), EDAC_ERROR(6) => 
        EDAC_ERROR(6), EDAC_ERROR(5) => EDAC_ERROR(5), 
        EDAC_ERROR(4) => EDAC_ERROR(4), EDAC_ERROR(3) => 
        EDAC_ERROR(3), EDAC_ERROR(2) => EDAC_ERROR(2), 
        EDAC_ERROR(1) => EDAC_ERROR(1), EDAC_ERROR(0) => 
        EDAC_ERROR(0), F_FM0_RDATA(31) => F_FM0_RDATA(31), 
        F_FM0_RDATA(30) => F_FM0_RDATA(30), F_FM0_RDATA(29) => 
        F_FM0_RDATA(29), F_FM0_RDATA(28) => F_FM0_RDATA(28), 
        F_FM0_RDATA(27) => F_FM0_RDATA(27), F_FM0_RDATA(26) => 
        F_FM0_RDATA(26), F_FM0_RDATA(25) => F_FM0_RDATA(25), 
        F_FM0_RDATA(24) => F_FM0_RDATA(24), F_FM0_RDATA(23) => 
        F_FM0_RDATA(23), F_FM0_RDATA(22) => F_FM0_RDATA(22), 
        F_FM0_RDATA(21) => F_FM0_RDATA(21), F_FM0_RDATA(20) => 
        F_FM0_RDATA(20), F_FM0_RDATA(19) => F_FM0_RDATA(19), 
        F_FM0_RDATA(18) => F_FM0_RDATA(18), F_FM0_RDATA(17) => 
        F_FM0_RDATA(17), F_FM0_RDATA(16) => F_FM0_RDATA(16), 
        F_FM0_RDATA(15) => F_FM0_RDATA(15), F_FM0_RDATA(14) => 
        F_FM0_RDATA(14), F_FM0_RDATA(13) => F_FM0_RDATA(13), 
        F_FM0_RDATA(12) => F_FM0_RDATA(12), F_FM0_RDATA(11) => 
        F_FM0_RDATA(11), F_FM0_RDATA(10) => F_FM0_RDATA(10), 
        F_FM0_RDATA(9) => F_FM0_RDATA(9), F_FM0_RDATA(8) => 
        F_FM0_RDATA(8), F_FM0_RDATA(7) => F_FM0_RDATA(7), 
        F_FM0_RDATA(6) => F_FM0_RDATA(6), F_FM0_RDATA(5) => 
        F_FM0_RDATA(5), F_FM0_RDATA(4) => F_FM0_RDATA(4), 
        F_FM0_RDATA(3) => F_FM0_RDATA(3), F_FM0_RDATA(2) => 
        F_FM0_RDATA(2), F_FM0_RDATA(1) => F_FM0_RDATA(1), 
        F_FM0_RDATA(0) => F_FM0_RDATA(0), F_FM0_READYOUT => 
        F_FM0_READYOUT, F_FM0_RESP => F_FM0_RESP, F_HM0_ADDR(31)
         => FIC_0_APB_M_PADDR(31), F_HM0_ADDR(30) => 
        FIC_0_APB_M_PADDR(30), F_HM0_ADDR(29) => 
        FIC_0_APB_M_PADDR(29), F_HM0_ADDR(28) => 
        FIC_0_APB_M_PADDR(28), F_HM0_ADDR(27) => 
        FIC_0_APB_M_PADDR(27), F_HM0_ADDR(26) => 
        FIC_0_APB_M_PADDR(26), F_HM0_ADDR(25) => 
        FIC_0_APB_M_PADDR(25), F_HM0_ADDR(24) => 
        FIC_0_APB_M_PADDR(24), F_HM0_ADDR(23) => 
        FIC_0_APB_M_PADDR(23), F_HM0_ADDR(22) => 
        FIC_0_APB_M_PADDR(22), F_HM0_ADDR(21) => 
        FIC_0_APB_M_PADDR(21), F_HM0_ADDR(20) => 
        FIC_0_APB_M_PADDR(20), F_HM0_ADDR(19) => 
        FIC_0_APB_M_PADDR(19), F_HM0_ADDR(18) => 
        FIC_0_APB_M_PADDR(18), F_HM0_ADDR(17) => 
        FIC_0_APB_M_PADDR(17), F_HM0_ADDR(16) => 
        FIC_0_APB_M_PADDR(16), F_HM0_ADDR(15) => STAMP_PADDRS(15), 
        F_HM0_ADDR(14) => STAMP_PADDRS(14), F_HM0_ADDR(13) => 
        STAMP_PADDRS(13), F_HM0_ADDR(12) => STAMP_PADDRS(12), 
        F_HM0_ADDR(11) => sb_sb_0_STAMP_PADDR(11), F_HM0_ADDR(10)
         => sb_sb_0_STAMP_PADDR(10), F_HM0_ADDR(9) => 
        sb_sb_0_STAMP_PADDR(9), F_HM0_ADDR(8) => 
        sb_sb_0_STAMP_PADDR(8), F_HM0_ADDR(7) => 
        sb_sb_0_STAMP_PADDR(7), F_HM0_ADDR(6) => 
        sb_sb_0_STAMP_PADDR(6), F_HM0_ADDR(5) => 
        sb_sb_0_STAMP_PADDR(5), F_HM0_ADDR(4) => 
        sb_sb_0_STAMP_PADDR(4), F_HM0_ADDR(3) => 
        sb_sb_0_STAMP_PADDR(3), F_HM0_ADDR(2) => 
        sb_sb_0_STAMP_PADDR(2), F_HM0_ADDR(1) => 
        sb_sb_0_STAMP_PADDR(1), F_HM0_ADDR(0) => 
        sb_sb_0_STAMP_PADDR(0), F_HM0_ENABLE => 
        sb_sb_0_STAMP_PENABLE, F_HM0_SEL => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, F_HM0_SIZE(1) => 
        F_HM0_SIZE(1), F_HM0_SIZE(0) => F_HM0_SIZE(0), 
        F_HM0_TRANS1 => F_HM0_TRANS1, F_HM0_WDATA(31) => 
        sb_sb_0_STAMP_PWDATA(31), F_HM0_WDATA(30) => 
        sb_sb_0_STAMP_PWDATA(30), F_HM0_WDATA(29) => 
        sb_sb_0_STAMP_PWDATA(29), F_HM0_WDATA(28) => 
        sb_sb_0_STAMP_PWDATA(28), F_HM0_WDATA(27) => 
        sb_sb_0_STAMP_PWDATA(27), F_HM0_WDATA(26) => 
        sb_sb_0_STAMP_PWDATA(26), F_HM0_WDATA(25) => 
        sb_sb_0_STAMP_PWDATA(25), F_HM0_WDATA(24) => 
        sb_sb_0_STAMP_PWDATA(24), F_HM0_WDATA(23) => 
        sb_sb_0_STAMP_PWDATA(23), F_HM0_WDATA(22) => 
        sb_sb_0_STAMP_PWDATA(22), F_HM0_WDATA(21) => 
        sb_sb_0_STAMP_PWDATA(21), F_HM0_WDATA(20) => 
        sb_sb_0_STAMP_PWDATA(20), F_HM0_WDATA(19) => 
        sb_sb_0_STAMP_PWDATA(19), F_HM0_WDATA(18) => 
        sb_sb_0_STAMP_PWDATA(18), F_HM0_WDATA(17) => 
        sb_sb_0_STAMP_PWDATA(17), F_HM0_WDATA(16) => 
        sb_sb_0_STAMP_PWDATA(16), F_HM0_WDATA(15) => 
        sb_sb_0_STAMP_PWDATA(15), F_HM0_WDATA(14) => 
        sb_sb_0_STAMP_PWDATA(14), F_HM0_WDATA(13) => 
        sb_sb_0_STAMP_PWDATA(13), F_HM0_WDATA(12) => 
        sb_sb_0_STAMP_PWDATA(12), F_HM0_WDATA(11) => 
        sb_sb_0_STAMP_PWDATA(11), F_HM0_WDATA(10) => 
        sb_sb_0_STAMP_PWDATA(10), F_HM0_WDATA(9) => 
        sb_sb_0_STAMP_PWDATA(9), F_HM0_WDATA(8) => 
        sb_sb_0_STAMP_PWDATA(8), F_HM0_WDATA(7) => 
        sb_sb_0_STAMP_PWDATA(7), F_HM0_WDATA(6) => 
        sb_sb_0_STAMP_PWDATA(6), F_HM0_WDATA(5) => 
        sb_sb_0_STAMP_PWDATA(5), F_HM0_WDATA(4) => 
        sb_sb_0_STAMP_PWDATA(4), F_HM0_WDATA(3) => 
        sb_sb_0_STAMP_PWDATA(3), F_HM0_WDATA(2) => 
        sb_sb_0_STAMP_PWDATA(2), F_HM0_WDATA(1) => 
        sb_sb_0_STAMP_PWDATA(1), F_HM0_WDATA(0) => 
        sb_sb_0_STAMP_PWDATA(0), F_HM0_WRITE => 
        sb_sb_0_STAMP_PWRITE, FAB_CHRGVBUS => FAB_CHRGVBUS, 
        FAB_DISCHRGVBUS => FAB_DISCHRGVBUS, FAB_DMPULLDOWN => 
        FAB_DMPULLDOWN, FAB_DPPULLDOWN => FAB_DPPULLDOWN, 
        FAB_DRVVBUS => FAB_DRVVBUS, FAB_IDPULLUP => FAB_IDPULLUP, 
        FAB_OPMODE(1) => FAB_OPMODE(1), FAB_OPMODE(0) => 
        FAB_OPMODE(0), FAB_SUSPENDM => FAB_SUSPENDM, FAB_TERMSEL
         => FAB_TERMSEL, FAB_TXVALID => FAB_TXVALID, 
        FAB_VCONTROL(3) => FAB_VCONTROL(3), FAB_VCONTROL(2) => 
        FAB_VCONTROL(2), FAB_VCONTROL(1) => FAB_VCONTROL(1), 
        FAB_VCONTROL(0) => FAB_VCONTROL(0), FAB_VCONTROLLOADM => 
        FAB_VCONTROLLOADM, FAB_XCVRSEL(1) => FAB_XCVRSEL(1), 
        FAB_XCVRSEL(0) => FAB_XCVRSEL(0), FAB_XDATAOUT(7) => 
        FAB_XDATAOUT(7), FAB_XDATAOUT(6) => FAB_XDATAOUT(6), 
        FAB_XDATAOUT(5) => FAB_XDATAOUT(5), FAB_XDATAOUT(4) => 
        FAB_XDATAOUT(4), FAB_XDATAOUT(3) => FAB_XDATAOUT(3), 
        FAB_XDATAOUT(2) => FAB_XDATAOUT(2), FAB_XDATAOUT(1) => 
        FAB_XDATAOUT(1), FAB_XDATAOUT(0) => FAB_XDATAOUT(0), 
        FACC_GLMUX_SEL => FACC_GLMUX_SEL, FIC32_0_MASTER(1) => 
        FIC32_0_MASTER(1), FIC32_0_MASTER(0) => FIC32_0_MASTER(0), 
        FIC32_1_MASTER(1) => FIC32_1_MASTER(1), FIC32_1_MASTER(0)
         => FIC32_1_MASTER(0), FPGA_RESET_N => MSS_RESET_N_M2F, 
        GTX_CLK => GTX_CLK, H2F_INTERRUPT(15) => 
        H2F_INTERRUPT(15), H2F_INTERRUPT(14) => H2F_INTERRUPT(14), 
        H2F_INTERRUPT(13) => H2F_INTERRUPT(13), H2F_INTERRUPT(12)
         => H2F_INTERRUPT(12), H2F_INTERRUPT(11) => 
        H2F_INTERRUPT(11), H2F_INTERRUPT(10) => H2F_INTERRUPT(10), 
        H2F_INTERRUPT(9) => H2F_INTERRUPT(9), H2F_INTERRUPT(8)
         => H2F_INTERRUPT(8), H2F_INTERRUPT(7) => 
        H2F_INTERRUPT(7), H2F_INTERRUPT(6) => H2F_INTERRUPT(6), 
        H2F_INTERRUPT(5) => H2F_INTERRUPT(5), H2F_INTERRUPT(4)
         => H2F_INTERRUPT(4), H2F_INTERRUPT(3) => 
        H2F_INTERRUPT(3), H2F_INTERRUPT(2) => H2F_INTERRUPT(2), 
        H2F_INTERRUPT(1) => H2F_INTERRUPT(1), H2F_INTERRUPT(0)
         => H2F_INTERRUPT(0), H2F_NMI => H2F_NMI, H2FCALIB => 
        H2FCALIB, I2C0_SCL_MGPIO31B_H2F_A => 
        I2C0_SCL_MGPIO31B_H2F_A, I2C0_SCL_MGPIO31B_H2F_B => 
        LED_HEARTBEAT_c, I2C0_SDA_MGPIO30B_H2F_A => 
        I2C0_SDA_MGPIO30B_H2F_A, I2C0_SDA_MGPIO30B_H2F_B => 
        LED_RECORDING_c, I2C1_SCL_MGPIO1A_H2F_A => 
        I2C1_SCL_MGPIO1A_H2F_A, I2C1_SCL_MGPIO1A_H2F_B => 
        I2C1_SCL_MGPIO1A_H2F_B, I2C1_SDA_MGPIO0A_H2F_A => 
        I2C1_SDA_MGPIO0A_H2F_A, I2C1_SDA_MGPIO0A_H2F_B => 
        I2C1_SDA_MGPIO0A_H2F_B, MDCF => MDCF, MDOENF => MDOENF, 
        MDOF => MDOF, MMUART0_CTS_MGPIO19B_H2F_A => 
        MMUART0_CTS_MGPIO19B_H2F_A, MMUART0_CTS_MGPIO19B_H2F_B
         => MMUART0_CTS_MGPIO19B_H2F_B, 
        MMUART0_DCD_MGPIO22B_H2F_A => MMUART0_DCD_MGPIO22B_H2F_A, 
        MMUART0_DCD_MGPIO22B_H2F_B => MMUART0_DCD_MGPIO22B_H2F_B, 
        MMUART0_DSR_MGPIO20B_H2F_A => MMUART0_DSR_MGPIO20B_H2F_A, 
        MMUART0_DSR_MGPIO20B_H2F_B => MMUART0_DSR_MGPIO20B_H2F_B, 
        MMUART0_DTR_MGPIO18B_H2F_A => MMUART0_DTR_MGPIO18B_H2F_A, 
        MMUART0_DTR_MGPIO18B_H2F_B => MMUART0_DTR_MGPIO18B_H2F_B, 
        MMUART0_RI_MGPIO21B_H2F_A => MMUART0_RI_MGPIO21B_H2F_A, 
        MMUART0_RI_MGPIO21B_H2F_B => MMUART0_RI_MGPIO21B_H2F_B, 
        MMUART0_RTS_MGPIO17B_H2F_A => MMUART0_RTS_MGPIO17B_H2F_A, 
        MMUART0_RTS_MGPIO17B_H2F_B => MMUART0_RTS_MGPIO17B_H2F_B, 
        MMUART0_RXD_MGPIO28B_H2F_A => MMUART0_RXD_MGPIO28B_H2F_A, 
        MMUART0_RXD_MGPIO28B_H2F_B => MMUART0_RXD_MGPIO28B_H2F_B, 
        MMUART0_SCK_MGPIO29B_H2F_A => MMUART0_SCK_MGPIO29B_H2F_A, 
        MMUART0_SCK_MGPIO29B_H2F_B => MMUART0_SCK_MGPIO29B_H2F_B, 
        MMUART0_TXD_MGPIO27B_H2F_A => MMUART0_TXD_MGPIO27B_H2F_A, 
        MMUART0_TXD_MGPIO27B_H2F_B => MMUART0_TXD_MGPIO27B_H2F_B, 
        MMUART1_DTR_MGPIO12B_H2F_A => MMUART1_DTR_MGPIO12B_H2F_A, 
        MMUART1_RTS_MGPIO11B_H2F_A => MMUART1_RTS_MGPIO11B_H2F_A, 
        MMUART1_RTS_MGPIO11B_H2F_B => MMUART1_RTS_MGPIO11B_H2F_B, 
        MMUART1_RXD_MGPIO26B_H2F_A => MMUART1_RXD_MGPIO26B_H2F_A, 
        MMUART1_RXD_MGPIO26B_H2F_B => MMUART1_RXD_MGPIO26B_H2F_B, 
        MMUART1_SCK_MGPIO25B_H2F_A => MMUART1_SCK_MGPIO25B_H2F_A, 
        MMUART1_SCK_MGPIO25B_H2F_B => MMUART1_SCK_MGPIO25B_H2F_B, 
        MMUART1_TXD_MGPIO24B_H2F_A => MMUART1_TXD_MGPIO24B_H2F_A, 
        MMUART1_TXD_MGPIO24B_H2F_B => MMUART1_TXD_MGPIO24B_H2F_B, 
        MPLL_LOCK => MPLL_LOCK, PER2_FABRIC_PADDR(15) => 
        FIC_2_APB_M_PADDR(15), PER2_FABRIC_PADDR(14) => 
        FIC_2_APB_M_PADDR(14), PER2_FABRIC_PADDR(13) => 
        FIC_2_APB_M_PADDR(13), PER2_FABRIC_PADDR(12) => 
        FIC_2_APB_M_PADDR(12), PER2_FABRIC_PADDR(11) => 
        FIC_2_APB_M_PADDR(11), PER2_FABRIC_PADDR(10) => 
        FIC_2_APB_M_PADDR(10), PER2_FABRIC_PADDR(9) => 
        FIC_2_APB_M_PADDR(9), PER2_FABRIC_PADDR(8) => 
        FIC_2_APB_M_PADDR(8), PER2_FABRIC_PADDR(7) => 
        FIC_2_APB_M_PADDR(7), PER2_FABRIC_PADDR(6) => 
        FIC_2_APB_M_PADDR(6), PER2_FABRIC_PADDR(5) => 
        FIC_2_APB_M_PADDR(5), PER2_FABRIC_PADDR(4) => 
        FIC_2_APB_M_PADDR(4), PER2_FABRIC_PADDR(3) => 
        FIC_2_APB_M_PADDR(3), PER2_FABRIC_PADDR(2) => 
        FIC_2_APB_M_PADDR(2), PER2_FABRIC_PENABLE => 
        FIC_2_APB_M_PENABLE, PER2_FABRIC_PSEL => FIC_2_APB_M_PSEL, 
        PER2_FABRIC_PWDATA(31) => FIC_2_APB_M_PWDATA(31), 
        PER2_FABRIC_PWDATA(30) => FIC_2_APB_M_PWDATA(30), 
        PER2_FABRIC_PWDATA(29) => FIC_2_APB_M_PWDATA(29), 
        PER2_FABRIC_PWDATA(28) => FIC_2_APB_M_PWDATA(28), 
        PER2_FABRIC_PWDATA(27) => FIC_2_APB_M_PWDATA(27), 
        PER2_FABRIC_PWDATA(26) => FIC_2_APB_M_PWDATA(26), 
        PER2_FABRIC_PWDATA(25) => FIC_2_APB_M_PWDATA(25), 
        PER2_FABRIC_PWDATA(24) => FIC_2_APB_M_PWDATA(24), 
        PER2_FABRIC_PWDATA(23) => FIC_2_APB_M_PWDATA(23), 
        PER2_FABRIC_PWDATA(22) => FIC_2_APB_M_PWDATA(22), 
        PER2_FABRIC_PWDATA(21) => FIC_2_APB_M_PWDATA(21), 
        PER2_FABRIC_PWDATA(20) => FIC_2_APB_M_PWDATA(20), 
        PER2_FABRIC_PWDATA(19) => FIC_2_APB_M_PWDATA(19), 
        PER2_FABRIC_PWDATA(18) => FIC_2_APB_M_PWDATA(18), 
        PER2_FABRIC_PWDATA(17) => FIC_2_APB_M_PWDATA(17), 
        PER2_FABRIC_PWDATA(16) => FIC_2_APB_M_PWDATA(16), 
        PER2_FABRIC_PWDATA(15) => FIC_2_APB_M_PWDATA(15), 
        PER2_FABRIC_PWDATA(14) => FIC_2_APB_M_PWDATA(14), 
        PER2_FABRIC_PWDATA(13) => FIC_2_APB_M_PWDATA(13), 
        PER2_FABRIC_PWDATA(12) => FIC_2_APB_M_PWDATA(12), 
        PER2_FABRIC_PWDATA(11) => FIC_2_APB_M_PWDATA(11), 
        PER2_FABRIC_PWDATA(10) => FIC_2_APB_M_PWDATA(10), 
        PER2_FABRIC_PWDATA(9) => FIC_2_APB_M_PWDATA(9), 
        PER2_FABRIC_PWDATA(8) => FIC_2_APB_M_PWDATA(8), 
        PER2_FABRIC_PWDATA(7) => FIC_2_APB_M_PWDATA(7), 
        PER2_FABRIC_PWDATA(6) => FIC_2_APB_M_PWDATA(6), 
        PER2_FABRIC_PWDATA(5) => FIC_2_APB_M_PWDATA(5), 
        PER2_FABRIC_PWDATA(4) => FIC_2_APB_M_PWDATA(4), 
        PER2_FABRIC_PWDATA(3) => FIC_2_APB_M_PWDATA(3), 
        PER2_FABRIC_PWDATA(2) => FIC_2_APB_M_PWDATA(2), 
        PER2_FABRIC_PWDATA(1) => FIC_2_APB_M_PWDATA(1), 
        PER2_FABRIC_PWDATA(0) => FIC_2_APB_M_PWDATA(0), 
        PER2_FABRIC_PWRITE => FIC_2_APB_M_PWRITE, RTC_MATCH => 
        RTC_MATCH, SLEEPDEEP => SLEEPDEEP, SLEEPHOLDACK => 
        SLEEPHOLDACK, SLEEPING => SLEEPING, SMBALERT_NO0 => 
        SMBALERT_NO0, SMBALERT_NO1 => SMBALERT_NO1, SMBSUS_NO0
         => SMBSUS_NO0, SMBSUS_NO1 => SMBSUS_NO1, SPI0_CLK_OUT
         => SPI0_CLK_OUT, SPI0_SDI_MGPIO5A_H2F_A => 
        SPI0_SDI_MGPIO5A_H2F_A, SPI0_SDI_MGPIO5A_H2F_B => 
        SPI0_SDI_MGPIO5A_H2F_B, SPI0_SDO_MGPIO6A_H2F_A => 
        SPI0_SDO_MGPIO6A_H2F_A, SPI0_SDO_MGPIO6A_H2F_B => 
        GPIO_6_M2F_c, SPI0_SS0_MGPIO7A_H2F_A => 
        SPI0_SS0_MGPIO7A_H2F_A, SPI0_SS0_MGPIO7A_H2F_B => 
        SPI0_SS0_MGPIO7A_H2F_B, SPI0_SS1_MGPIO8A_H2F_A => 
        SPI0_SS1_MGPIO8A_H2F_A, SPI0_SS1_MGPIO8A_H2F_B => 
        SPI0_SS1_MGPIO8A_H2F_B, SPI0_SS2_MGPIO9A_H2F_A => 
        SPI0_SS2_MGPIO9A_H2F_A, SPI0_SS2_MGPIO9A_H2F_B => 
        SPI0_SS2_MGPIO9A_H2F_B, SPI0_SS3_MGPIO10A_H2F_A => 
        SPI0_SS3_MGPIO10A_H2F_A, SPI0_SS3_MGPIO10A_H2F_B => 
        SPI0_SS3_MGPIO10A_H2F_B, SPI0_SS4_MGPIO19A_H2F_A => 
        SPI0_SS4_MGPIO19A_H2F_A, SPI0_SS5_MGPIO20A_H2F_A => 
        SPI0_SS5_MGPIO20A_H2F_A, SPI0_SS6_MGPIO21A_H2F_A => 
        SPI0_SS6_MGPIO21A_H2F_A, SPI0_SS7_MGPIO22A_H2F_A => 
        SPI0_SS7_MGPIO22A_H2F_A, SPI1_CLK_OUT => SPI1_CLK_OUT, 
        SPI1_SDI_MGPIO11A_H2F_A => SPI1_SDI_MGPIO11A_H2F_A, 
        SPI1_SDI_MGPIO11A_H2F_B => SPI1_SDI_MGPIO11A_H2F_B, 
        SPI1_SDO_MGPIO12A_H2F_A => SPI1_SDO_MGPIO12A_H2F_A, 
        SPI1_SDO_MGPIO12A_H2F_B => SPI1_SDO_MGPIO12A_H2F_B, 
        SPI1_SS0_MGPIO13A_H2F_A => SPI1_SS0_MGPIO13A_H2F_A, 
        SPI1_SS0_MGPIO13A_H2F_B => SPI1_SS0_MGPIO13A_H2F_B, 
        SPI1_SS1_MGPIO14A_H2F_A => SPI1_SS1_MGPIO14A_H2F_A, 
        SPI1_SS1_MGPIO14A_H2F_B => SPI1_SS1_MGPIO14A_H2F_B, 
        SPI1_SS2_MGPIO15A_H2F_A => SPI1_SS2_MGPIO15A_H2F_A, 
        SPI1_SS2_MGPIO15A_H2F_B => SPI1_SS2_MGPIO15A_H2F_B, 
        SPI1_SS3_MGPIO16A_H2F_A => SPI1_SS3_MGPIO16A_H2F_A, 
        SPI1_SS3_MGPIO16A_H2F_B => SPI1_SS3_MGPIO16A_H2F_B, 
        SPI1_SS4_MGPIO17A_H2F_A => SPI1_SS4_MGPIO17A_H2F_A, 
        SPI1_SS5_MGPIO18A_H2F_A => SPI1_SS5_MGPIO18A_H2F_A, 
        SPI1_SS6_MGPIO23A_H2F_A => SPI1_SS6_MGPIO23A_H2F_A, 
        SPI1_SS7_MGPIO24A_H2F_A => SPI1_SS7_MGPIO24A_H2F_A, 
        TCGF(9) => TCGF(9), TCGF(8) => TCGF(8), TCGF(7) => 
        TCGF(7), TCGF(6) => TCGF(6), TCGF(5) => TCGF(5), TCGF(4)
         => TCGF(4), TCGF(3) => TCGF(3), TCGF(2) => TCGF(2), 
        TCGF(1) => TCGF(1), TCGF(0) => TCGF(0), TRACECLK => 
        TRACECLK, TRACEDATA(3) => TRACEDATA(3), TRACEDATA(2) => 
        TRACEDATA(2), TRACEDATA(1) => TRACEDATA(1), TRACEDATA(0)
         => TRACEDATA(0), TX_CLK => TX_CLK, TX_ENF => TX_ENF, 
        TX_ERRF => TX_ERRF, TXCTL_EN_RIF => TXCTL_EN_RIF, 
        TXD_RIF(3) => TXD_RIF(3), TXD_RIF(2) => TXD_RIF(2), 
        TXD_RIF(1) => TXD_RIF(1), TXD_RIF(0) => TXD_RIF(0), 
        TXDF(7) => TXDF(7), TXDF(6) => TXDF(6), TXDF(5) => 
        TXDF(5), TXDF(4) => TXDF(4), TXDF(3) => TXDF(3), TXDF(2)
         => TXDF(2), TXDF(1) => TXDF(1), TXDF(0) => TXDF(0), TXEV
         => TXEV, WDOGTIMEOUT => WDOGTIMEOUT, 
        F_ARREADY_HREADYOUT1 => F_ARREADY_HREADYOUT1, 
        F_AWREADY_HREADYOUT0 => F_AWREADY_HREADYOUT0, F_BID(3)
         => F_BID(3), F_BID(2) => F_BID(2), F_BID(1) => F_BID(1), 
        F_BID(0) => F_BID(0), F_BRESP_HRESP0(1) => 
        F_BRESP_HRESP0(1), F_BRESP_HRESP0(0) => F_BRESP_HRESP0(0), 
        F_BVALID => F_BVALID, F_RDATA_HRDATA01(63) => 
        F_RDATA_HRDATA01(63), F_RDATA_HRDATA01(62) => 
        F_RDATA_HRDATA01(62), F_RDATA_HRDATA01(61) => 
        F_RDATA_HRDATA01(61), F_RDATA_HRDATA01(60) => 
        F_RDATA_HRDATA01(60), F_RDATA_HRDATA01(59) => 
        F_RDATA_HRDATA01(59), F_RDATA_HRDATA01(58) => 
        F_RDATA_HRDATA01(58), F_RDATA_HRDATA01(57) => 
        F_RDATA_HRDATA01(57), F_RDATA_HRDATA01(56) => 
        F_RDATA_HRDATA01(56), F_RDATA_HRDATA01(55) => 
        F_RDATA_HRDATA01(55), F_RDATA_HRDATA01(54) => 
        F_RDATA_HRDATA01(54), F_RDATA_HRDATA01(53) => 
        F_RDATA_HRDATA01(53), F_RDATA_HRDATA01(52) => 
        F_RDATA_HRDATA01(52), F_RDATA_HRDATA01(51) => 
        F_RDATA_HRDATA01(51), F_RDATA_HRDATA01(50) => 
        F_RDATA_HRDATA01(50), F_RDATA_HRDATA01(49) => 
        F_RDATA_HRDATA01(49), F_RDATA_HRDATA01(48) => 
        F_RDATA_HRDATA01(48), F_RDATA_HRDATA01(47) => 
        F_RDATA_HRDATA01(47), F_RDATA_HRDATA01(46) => 
        F_RDATA_HRDATA01(46), F_RDATA_HRDATA01(45) => 
        F_RDATA_HRDATA01(45), F_RDATA_HRDATA01(44) => 
        F_RDATA_HRDATA01(44), F_RDATA_HRDATA01(43) => 
        F_RDATA_HRDATA01(43), F_RDATA_HRDATA01(42) => 
        F_RDATA_HRDATA01(42), F_RDATA_HRDATA01(41) => 
        F_RDATA_HRDATA01(41), F_RDATA_HRDATA01(40) => 
        F_RDATA_HRDATA01(40), F_RDATA_HRDATA01(39) => 
        F_RDATA_HRDATA01(39), F_RDATA_HRDATA01(38) => 
        F_RDATA_HRDATA01(38), F_RDATA_HRDATA01(37) => 
        F_RDATA_HRDATA01(37), F_RDATA_HRDATA01(36) => 
        F_RDATA_HRDATA01(36), F_RDATA_HRDATA01(35) => 
        F_RDATA_HRDATA01(35), F_RDATA_HRDATA01(34) => 
        F_RDATA_HRDATA01(34), F_RDATA_HRDATA01(33) => 
        F_RDATA_HRDATA01(33), F_RDATA_HRDATA01(32) => 
        F_RDATA_HRDATA01(32), F_RDATA_HRDATA01(31) => 
        F_RDATA_HRDATA01(31), F_RDATA_HRDATA01(30) => 
        F_RDATA_HRDATA01(30), F_RDATA_HRDATA01(29) => 
        F_RDATA_HRDATA01(29), F_RDATA_HRDATA01(28) => 
        F_RDATA_HRDATA01(28), F_RDATA_HRDATA01(27) => 
        F_RDATA_HRDATA01(27), F_RDATA_HRDATA01(26) => 
        F_RDATA_HRDATA01(26), F_RDATA_HRDATA01(25) => 
        F_RDATA_HRDATA01(25), F_RDATA_HRDATA01(24) => 
        F_RDATA_HRDATA01(24), F_RDATA_HRDATA01(23) => 
        F_RDATA_HRDATA01(23), F_RDATA_HRDATA01(22) => 
        F_RDATA_HRDATA01(22), F_RDATA_HRDATA01(21) => 
        F_RDATA_HRDATA01(21), F_RDATA_HRDATA01(20) => 
        F_RDATA_HRDATA01(20), F_RDATA_HRDATA01(19) => 
        F_RDATA_HRDATA01(19), F_RDATA_HRDATA01(18) => 
        F_RDATA_HRDATA01(18), F_RDATA_HRDATA01(17) => 
        F_RDATA_HRDATA01(17), F_RDATA_HRDATA01(16) => 
        F_RDATA_HRDATA01(16), F_RDATA_HRDATA01(15) => 
        F_RDATA_HRDATA01(15), F_RDATA_HRDATA01(14) => 
        F_RDATA_HRDATA01(14), F_RDATA_HRDATA01(13) => 
        F_RDATA_HRDATA01(13), F_RDATA_HRDATA01(12) => 
        F_RDATA_HRDATA01(12), F_RDATA_HRDATA01(11) => 
        F_RDATA_HRDATA01(11), F_RDATA_HRDATA01(10) => 
        F_RDATA_HRDATA01(10), F_RDATA_HRDATA01(9) => 
        F_RDATA_HRDATA01(9), F_RDATA_HRDATA01(8) => 
        F_RDATA_HRDATA01(8), F_RDATA_HRDATA01(7) => 
        F_RDATA_HRDATA01(7), F_RDATA_HRDATA01(6) => 
        F_RDATA_HRDATA01(6), F_RDATA_HRDATA01(5) => 
        F_RDATA_HRDATA01(5), F_RDATA_HRDATA01(4) => 
        F_RDATA_HRDATA01(4), F_RDATA_HRDATA01(3) => 
        F_RDATA_HRDATA01(3), F_RDATA_HRDATA01(2) => 
        F_RDATA_HRDATA01(2), F_RDATA_HRDATA01(1) => 
        F_RDATA_HRDATA01(1), F_RDATA_HRDATA01(0) => 
        F_RDATA_HRDATA01(0), F_RID(3) => F_RID(3), F_RID(2) => 
        F_RID(2), F_RID(1) => F_RID(1), F_RID(0) => F_RID(0), 
        F_RLAST => F_RLAST, F_RRESP_HRESP1(1) => 
        F_RRESP_HRESP1(1), F_RRESP_HRESP1(0) => F_RRESP_HRESP1(0), 
        F_RVALID => F_RVALID, F_WREADY => F_WREADY, 
        MDDR_FABRIC_PRDATA(15) => MDDR_FABRIC_PRDATA(15), 
        MDDR_FABRIC_PRDATA(14) => MDDR_FABRIC_PRDATA(14), 
        MDDR_FABRIC_PRDATA(13) => MDDR_FABRIC_PRDATA(13), 
        MDDR_FABRIC_PRDATA(12) => MDDR_FABRIC_PRDATA(12), 
        MDDR_FABRIC_PRDATA(11) => MDDR_FABRIC_PRDATA(11), 
        MDDR_FABRIC_PRDATA(10) => MDDR_FABRIC_PRDATA(10), 
        MDDR_FABRIC_PRDATA(9) => MDDR_FABRIC_PRDATA(9), 
        MDDR_FABRIC_PRDATA(8) => MDDR_FABRIC_PRDATA(8), 
        MDDR_FABRIC_PRDATA(7) => MDDR_FABRIC_PRDATA(7), 
        MDDR_FABRIC_PRDATA(6) => MDDR_FABRIC_PRDATA(6), 
        MDDR_FABRIC_PRDATA(5) => MDDR_FABRIC_PRDATA(5), 
        MDDR_FABRIC_PRDATA(4) => MDDR_FABRIC_PRDATA(4), 
        MDDR_FABRIC_PRDATA(3) => MDDR_FABRIC_PRDATA(3), 
        MDDR_FABRIC_PRDATA(2) => MDDR_FABRIC_PRDATA(2), 
        MDDR_FABRIC_PRDATA(1) => MDDR_FABRIC_PRDATA(1), 
        MDDR_FABRIC_PRDATA(0) => MDDR_FABRIC_PRDATA(0), 
        MDDR_FABRIC_PREADY => MDDR_FABRIC_PREADY, 
        MDDR_FABRIC_PSLVERR => MDDR_FABRIC_PSLVERR, 
        CAN_RXBUS_F2H_SCP => \VCC\, CAN_TX_EBL_F2H_SCP => \VCC\, 
        CAN_TXBUS_F2H_SCP => \VCC\, COLF => \VCC\, CRSF => \VCC\, 
        F2_DMAREADY(1) => \VCC\, F2_DMAREADY(0) => \VCC\, 
        F2H_INTERRUPT(15) => \GND\, F2H_INTERRUPT(14) => \GND\, 
        F2H_INTERRUPT(13) => \GND\, F2H_INTERRUPT(12) => \GND\, 
        F2H_INTERRUPT(11) => \GND\, F2H_INTERRUPT(10) => \GND\, 
        F2H_INTERRUPT(9) => \GND\, F2H_INTERRUPT(8) => \GND\, 
        F2H_INTERRUPT(7) => \GND\, F2H_INTERRUPT(6) => \GND\, 
        F2H_INTERRUPT(5) => \GND\, F2H_INTERRUPT(4) => \GND\, 
        F2H_INTERRUPT(3) => \GND\, F2H_INTERRUPT(2) => \GND\, 
        F2H_INTERRUPT(1) => \GND\, F2H_INTERRUPT(0) => 
        dataReady_0, F2HCALIB => \VCC\, F_DMAREADY(1) => \VCC\, 
        F_DMAREADY(0) => \VCC\, F_FM0_ADDR(31) => \GND\, 
        F_FM0_ADDR(30) => \GND\, F_FM0_ADDR(29) => \GND\, 
        F_FM0_ADDR(28) => \GND\, F_FM0_ADDR(27) => \GND\, 
        F_FM0_ADDR(26) => \GND\, F_FM0_ADDR(25) => \GND\, 
        F_FM0_ADDR(24) => \GND\, F_FM0_ADDR(23) => \GND\, 
        F_FM0_ADDR(22) => \GND\, F_FM0_ADDR(21) => \GND\, 
        F_FM0_ADDR(20) => \GND\, F_FM0_ADDR(19) => \GND\, 
        F_FM0_ADDR(18) => \GND\, F_FM0_ADDR(17) => \GND\, 
        F_FM0_ADDR(16) => \GND\, F_FM0_ADDR(15) => \GND\, 
        F_FM0_ADDR(14) => \GND\, F_FM0_ADDR(13) => \GND\, 
        F_FM0_ADDR(12) => \GND\, F_FM0_ADDR(11) => \GND\, 
        F_FM0_ADDR(10) => \GND\, F_FM0_ADDR(9) => \GND\, 
        F_FM0_ADDR(8) => \GND\, F_FM0_ADDR(7) => \GND\, 
        F_FM0_ADDR(6) => \GND\, F_FM0_ADDR(5) => \GND\, 
        F_FM0_ADDR(4) => \GND\, F_FM0_ADDR(3) => \GND\, 
        F_FM0_ADDR(2) => \GND\, F_FM0_ADDR(1) => \GND\, 
        F_FM0_ADDR(0) => \GND\, F_FM0_ENABLE => \GND\, 
        F_FM0_MASTLOCK => \GND\, F_FM0_READY => \VCC\, F_FM0_SEL
         => \GND\, F_FM0_SIZE(1) => \GND\, F_FM0_SIZE(0) => \GND\, 
        F_FM0_TRANS1 => \GND\, F_FM0_WDATA(31) => \GND\, 
        F_FM0_WDATA(30) => \GND\, F_FM0_WDATA(29) => \GND\, 
        F_FM0_WDATA(28) => \GND\, F_FM0_WDATA(27) => \GND\, 
        F_FM0_WDATA(26) => \GND\, F_FM0_WDATA(25) => \GND\, 
        F_FM0_WDATA(24) => \GND\, F_FM0_WDATA(23) => \GND\, 
        F_FM0_WDATA(22) => \GND\, F_FM0_WDATA(21) => \GND\, 
        F_FM0_WDATA(20) => \GND\, F_FM0_WDATA(19) => \GND\, 
        F_FM0_WDATA(18) => \GND\, F_FM0_WDATA(17) => \GND\, 
        F_FM0_WDATA(16) => \GND\, F_FM0_WDATA(15) => \GND\, 
        F_FM0_WDATA(14) => \GND\, F_FM0_WDATA(13) => \GND\, 
        F_FM0_WDATA(12) => \GND\, F_FM0_WDATA(11) => \GND\, 
        F_FM0_WDATA(10) => \GND\, F_FM0_WDATA(9) => \GND\, 
        F_FM0_WDATA(8) => \GND\, F_FM0_WDATA(7) => \GND\, 
        F_FM0_WDATA(6) => \GND\, F_FM0_WDATA(5) => \GND\, 
        F_FM0_WDATA(4) => \GND\, F_FM0_WDATA(3) => \GND\, 
        F_FM0_WDATA(2) => \GND\, F_FM0_WDATA(1) => \GND\, 
        F_FM0_WDATA(0) => \GND\, F_FM0_WRITE => \GND\, 
        F_HM0_RDATA(31) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31), 
        F_HM0_RDATA(30) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30), 
        F_HM0_RDATA(29) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29), 
        F_HM0_RDATA(28) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28), 
        F_HM0_RDATA(27) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27), 
        F_HM0_RDATA(26) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26), 
        F_HM0_RDATA(25) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25), 
        F_HM0_RDATA(24) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24), 
        F_HM0_RDATA(23) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23), 
        F_HM0_RDATA(22) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22), 
        F_HM0_RDATA(21) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21), 
        F_HM0_RDATA(20) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20), 
        F_HM0_RDATA(19) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19), 
        F_HM0_RDATA(18) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18), 
        F_HM0_RDATA(17) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17), 
        F_HM0_RDATA(16) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16), 
        F_HM0_RDATA(15) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15), 
        F_HM0_RDATA(14) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14), 
        F_HM0_RDATA(13) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13), 
        F_HM0_RDATA(12) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12), 
        F_HM0_RDATA(11) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11), 
        F_HM0_RDATA(10) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10), 
        F_HM0_RDATA(9) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9), 
        F_HM0_RDATA(8) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8), 
        F_HM0_RDATA(7) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(7), 
        F_HM0_RDATA(6) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(6), 
        F_HM0_RDATA(5) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(5), 
        F_HM0_RDATA(4) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(4), 
        F_HM0_RDATA(3) => PRDATA_N_5_i, F_HM0_RDATA(2) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(2), 
        F_HM0_RDATA(1) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(1), 
        F_HM0_RDATA(0) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(0), F_HM0_READY
         => PREADY_N_7, F_HM0_RESP => \GND\, FAB_AVALID => \VCC\, 
        FAB_HOSTDISCON => \VCC\, FAB_IDDIG => \VCC\, 
        FAB_LINESTATE(1) => \VCC\, FAB_LINESTATE(0) => \VCC\, 
        FAB_M3_RESET_N => \VCC\, FAB_PLL_LOCK => FIC_0_LOCK, 
        FAB_RXACTIVE => \VCC\, FAB_RXERROR => \VCC\, FAB_RXVALID
         => \VCC\, FAB_RXVALIDH => \GND\, FAB_SESSEND => \VCC\, 
        FAB_TXREADY => \VCC\, FAB_VBUSVALID => \VCC\, 
        FAB_VSTATUS(7) => \VCC\, FAB_VSTATUS(6) => \VCC\, 
        FAB_VSTATUS(5) => \VCC\, FAB_VSTATUS(4) => \VCC\, 
        FAB_VSTATUS(3) => \VCC\, FAB_VSTATUS(2) => \VCC\, 
        FAB_VSTATUS(1) => \VCC\, FAB_VSTATUS(0) => \VCC\, 
        FAB_XDATAIN(7) => \VCC\, FAB_XDATAIN(6) => \VCC\, 
        FAB_XDATAIN(5) => \VCC\, FAB_XDATAIN(4) => \VCC\, 
        FAB_XDATAIN(3) => \VCC\, FAB_XDATAIN(2) => \VCC\, 
        FAB_XDATAIN(1) => \VCC\, FAB_XDATAIN(0) => \VCC\, 
        GTX_CLKPF => \VCC\, I2C0_BCLK => \VCC\, I2C0_SCL_F2H_SCP
         => \VCC\, I2C0_SDA_F2H_SCP => \VCC\, I2C1_BCLK => \VCC\, 
        I2C1_SCL_F2H_SCP => \VCC\, I2C1_SDA_F2H_SCP => \VCC\, 
        MDIF => \VCC\, MGPIO0A_F2H_GPIN => RXSM_LO_c, 
        MGPIO10A_F2H_GPIN => \VCC\, MGPIO11A_F2H_GPIN => \VCC\, 
        MGPIO11B_F2H_GPIN => \VCC\, MGPIO12A_F2H_GPIN => \VCC\, 
        MGPIO13A_F2H_GPIN => \VCC\, MGPIO14A_F2H_GPIN => \VCC\, 
        MGPIO15A_F2H_GPIN => \VCC\, MGPIO16A_F2H_GPIN => \VCC\, 
        MGPIO17B_F2H_GPIN => \VCC\, MGPIO18B_F2H_GPIN => \VCC\, 
        MGPIO19B_F2H_GPIN => \VCC\, MGPIO1A_F2H_GPIN => 
        RXSM_SOE_c, MGPIO20B_F2H_GPIN => \VCC\, MGPIO21B_F2H_GPIN
         => \VCC\, MGPIO22B_F2H_GPIN => \VCC\, MGPIO24B_F2H_GPIN
         => \VCC\, MGPIO25B_F2H_GPIN => \VCC\, MGPIO26B_F2H_GPIN
         => \VCC\, MGPIO27B_F2H_GPIN => \VCC\, MGPIO28B_F2H_GPIN
         => \VCC\, MGPIO29B_F2H_GPIN => \VCC\, MGPIO2A_F2H_GPIN
         => RXSM_SODS_c, MGPIO30B_F2H_GPIN => \VCC\, 
        MGPIO31B_F2H_GPIN => \VCC\, MGPIO3A_F2H_GPIN => \VCC\, 
        MGPIO4A_F2H_GPIN => \VCC\, MGPIO5A_F2H_GPIN => \VCC\, 
        MGPIO6A_F2H_GPIN => \VCC\, MGPIO7A_F2H_GPIN => \VCC\, 
        MGPIO8A_F2H_GPIN => \VCC\, MGPIO9A_F2H_GPIN => \VCC\, 
        MMUART0_CTS_F2H_SCP => \VCC\, MMUART0_DCD_F2H_SCP => 
        \VCC\, MMUART0_DSR_F2H_SCP => \VCC\, MMUART0_DTR_F2H_SCP
         => \VCC\, MMUART0_RI_F2H_SCP => \VCC\, 
        MMUART0_RTS_F2H_SCP => \VCC\, MMUART0_RXD_F2H_SCP => 
        \VCC\, MMUART0_SCK_F2H_SCP => \VCC\, MMUART0_TXD_F2H_SCP
         => \VCC\, MMUART1_CTS_F2H_SCP => \VCC\, 
        MMUART1_DCD_F2H_SCP => \VCC\, MMUART1_DSR_F2H_SCP => 
        \VCC\, MMUART1_RI_F2H_SCP => \VCC\, MMUART1_RTS_F2H_SCP
         => \VCC\, MMUART1_RXD_F2H_SCP => \VCC\, 
        MMUART1_SCK_F2H_SCP => \VCC\, MMUART1_TXD_F2H_SCP => 
        \VCC\, PER2_FABRIC_PRDATA(31) => \GND\, 
        PER2_FABRIC_PRDATA(30) => \GND\, PER2_FABRIC_PRDATA(29)
         => \GND\, PER2_FABRIC_PRDATA(28) => \GND\, 
        PER2_FABRIC_PRDATA(27) => \GND\, PER2_FABRIC_PRDATA(26)
         => \GND\, PER2_FABRIC_PRDATA(25) => \GND\, 
        PER2_FABRIC_PRDATA(24) => \GND\, PER2_FABRIC_PRDATA(23)
         => \GND\, PER2_FABRIC_PRDATA(22) => \GND\, 
        PER2_FABRIC_PRDATA(21) => \GND\, PER2_FABRIC_PRDATA(20)
         => \GND\, PER2_FABRIC_PRDATA(19) => \GND\, 
        PER2_FABRIC_PRDATA(18) => \GND\, PER2_FABRIC_PRDATA(17)
         => \GND\, PER2_FABRIC_PRDATA(16) => \GND\, 
        PER2_FABRIC_PRDATA(15) => \GND\, PER2_FABRIC_PRDATA(14)
         => \GND\, PER2_FABRIC_PRDATA(13) => \GND\, 
        PER2_FABRIC_PRDATA(12) => \GND\, PER2_FABRIC_PRDATA(11)
         => \GND\, PER2_FABRIC_PRDATA(10) => \GND\, 
        PER2_FABRIC_PRDATA(9) => \GND\, PER2_FABRIC_PRDATA(8) => 
        \GND\, PER2_FABRIC_PRDATA(7) => \GND\, 
        PER2_FABRIC_PRDATA(6) => \GND\, PER2_FABRIC_PRDATA(5) => 
        \GND\, PER2_FABRIC_PRDATA(4) => \GND\, 
        PER2_FABRIC_PRDATA(3) => \GND\, PER2_FABRIC_PRDATA(2) => 
        \GND\, PER2_FABRIC_PRDATA(1) => \GND\, 
        PER2_FABRIC_PRDATA(0) => \GND\, PER2_FABRIC_PREADY => 
        \VCC\, PER2_FABRIC_PSLVERR => \GND\, RCGF(9) => \VCC\, 
        RCGF(8) => \VCC\, RCGF(7) => \VCC\, RCGF(6) => \VCC\, 
        RCGF(5) => \VCC\, RCGF(4) => \VCC\, RCGF(3) => \VCC\, 
        RCGF(2) => \VCC\, RCGF(1) => \VCC\, RCGF(0) => \VCC\, 
        RX_CLKPF => \VCC\, RX_DVF => \VCC\, RX_ERRF => \VCC\, 
        RX_EV => \VCC\, RXDF(7) => \VCC\, RXDF(6) => \VCC\, 
        RXDF(5) => \VCC\, RXDF(4) => \VCC\, RXDF(3) => \VCC\, 
        RXDF(2) => \VCC\, RXDF(1) => \VCC\, RXDF(0) => \VCC\, 
        SLEEPHOLDREQ => \GND\, SMBALERT_NI0 => \VCC\, 
        SMBALERT_NI1 => \VCC\, SMBSUS_NI0 => \VCC\, SMBSUS_NI1
         => \VCC\, SPI0_CLK_IN => \VCC\, SPI0_SDI_F2H_SCP => 
        \VCC\, SPI0_SDO_F2H_SCP => \VCC\, SPI0_SS0_F2H_SCP => 
        \VCC\, SPI0_SS1_F2H_SCP => \VCC\, SPI0_SS2_F2H_SCP => 
        \VCC\, SPI0_SS3_F2H_SCP => \VCC\, SPI1_CLK_IN => \VCC\, 
        SPI1_SDI_F2H_SCP => \VCC\, SPI1_SDO_F2H_SCP => \VCC\, 
        SPI1_SS0_F2H_SCP => \VCC\, SPI1_SS1_F2H_SCP => \VCC\, 
        SPI1_SS2_F2H_SCP => \VCC\, SPI1_SS3_F2H_SCP => \VCC\, 
        TX_CLKPF => \VCC\, USER_MSS_GPIO_RESET_N => \VCC\, 
        USER_MSS_RESET_N => \VCC\, XCLK_FAB => \VCC\, CLK_BASE
         => sb_sb_0_FIC_0_CLK, CLK_MDDR_APB => \VCC\, 
        F_ARADDR_HADDR1(31) => \VCC\, F_ARADDR_HADDR1(30) => 
        \VCC\, F_ARADDR_HADDR1(29) => \VCC\, F_ARADDR_HADDR1(28)
         => \VCC\, F_ARADDR_HADDR1(27) => \VCC\, 
        F_ARADDR_HADDR1(26) => \VCC\, F_ARADDR_HADDR1(25) => 
        \VCC\, F_ARADDR_HADDR1(24) => \VCC\, F_ARADDR_HADDR1(23)
         => \VCC\, F_ARADDR_HADDR1(22) => \VCC\, 
        F_ARADDR_HADDR1(21) => \VCC\, F_ARADDR_HADDR1(20) => 
        \VCC\, F_ARADDR_HADDR1(19) => \VCC\, F_ARADDR_HADDR1(18)
         => \VCC\, F_ARADDR_HADDR1(17) => \VCC\, 
        F_ARADDR_HADDR1(16) => \VCC\, F_ARADDR_HADDR1(15) => 
        \VCC\, F_ARADDR_HADDR1(14) => \VCC\, F_ARADDR_HADDR1(13)
         => \VCC\, F_ARADDR_HADDR1(12) => \VCC\, 
        F_ARADDR_HADDR1(11) => \VCC\, F_ARADDR_HADDR1(10) => 
        \VCC\, F_ARADDR_HADDR1(9) => \VCC\, F_ARADDR_HADDR1(8)
         => \VCC\, F_ARADDR_HADDR1(7) => \VCC\, 
        F_ARADDR_HADDR1(6) => \VCC\, F_ARADDR_HADDR1(5) => \VCC\, 
        F_ARADDR_HADDR1(4) => \VCC\, F_ARADDR_HADDR1(3) => \VCC\, 
        F_ARADDR_HADDR1(2) => \VCC\, F_ARADDR_HADDR1(1) => \VCC\, 
        F_ARADDR_HADDR1(0) => \VCC\, F_ARBURST_HTRANS1(1) => 
        \GND\, F_ARBURST_HTRANS1(0) => \GND\, F_ARID_HSEL1(3) => 
        \GND\, F_ARID_HSEL1(2) => \GND\, F_ARID_HSEL1(1) => \GND\, 
        F_ARID_HSEL1(0) => \GND\, F_ARLEN_HBURST1(3) => \GND\, 
        F_ARLEN_HBURST1(2) => \GND\, F_ARLEN_HBURST1(1) => \GND\, 
        F_ARLEN_HBURST1(0) => \GND\, F_ARLOCK_HMASTLOCK1(1) => 
        \GND\, F_ARLOCK_HMASTLOCK1(0) => \GND\, 
        F_ARSIZE_HSIZE1(1) => \GND\, F_ARSIZE_HSIZE1(0) => \GND\, 
        F_ARVALID_HWRITE1 => \GND\, F_AWADDR_HADDR0(31) => \VCC\, 
        F_AWADDR_HADDR0(30) => \VCC\, F_AWADDR_HADDR0(29) => 
        \VCC\, F_AWADDR_HADDR0(28) => \VCC\, F_AWADDR_HADDR0(27)
         => \VCC\, F_AWADDR_HADDR0(26) => \VCC\, 
        F_AWADDR_HADDR0(25) => \VCC\, F_AWADDR_HADDR0(24) => 
        \VCC\, F_AWADDR_HADDR0(23) => \VCC\, F_AWADDR_HADDR0(22)
         => \VCC\, F_AWADDR_HADDR0(21) => \VCC\, 
        F_AWADDR_HADDR0(20) => \VCC\, F_AWADDR_HADDR0(19) => 
        \VCC\, F_AWADDR_HADDR0(18) => \VCC\, F_AWADDR_HADDR0(17)
         => \VCC\, F_AWADDR_HADDR0(16) => \VCC\, 
        F_AWADDR_HADDR0(15) => \VCC\, F_AWADDR_HADDR0(14) => 
        \VCC\, F_AWADDR_HADDR0(13) => \VCC\, F_AWADDR_HADDR0(12)
         => \VCC\, F_AWADDR_HADDR0(11) => \VCC\, 
        F_AWADDR_HADDR0(10) => \VCC\, F_AWADDR_HADDR0(9) => \VCC\, 
        F_AWADDR_HADDR0(8) => \VCC\, F_AWADDR_HADDR0(7) => \VCC\, 
        F_AWADDR_HADDR0(6) => \VCC\, F_AWADDR_HADDR0(5) => \VCC\, 
        F_AWADDR_HADDR0(4) => \VCC\, F_AWADDR_HADDR0(3) => \VCC\, 
        F_AWADDR_HADDR0(2) => \VCC\, F_AWADDR_HADDR0(1) => \VCC\, 
        F_AWADDR_HADDR0(0) => \VCC\, F_AWBURST_HTRANS0(1) => 
        \GND\, F_AWBURST_HTRANS0(0) => \GND\, F_AWID_HSEL0(3) => 
        \GND\, F_AWID_HSEL0(2) => \GND\, F_AWID_HSEL0(1) => \GND\, 
        F_AWID_HSEL0(0) => \GND\, F_AWLEN_HBURST0(3) => \GND\, 
        F_AWLEN_HBURST0(2) => \GND\, F_AWLEN_HBURST0(1) => \GND\, 
        F_AWLEN_HBURST0(0) => \GND\, F_AWLOCK_HMASTLOCK0(1) => 
        \GND\, F_AWLOCK_HMASTLOCK0(0) => \GND\, 
        F_AWSIZE_HSIZE0(1) => \GND\, F_AWSIZE_HSIZE0(0) => \GND\, 
        F_AWVALID_HWRITE0 => \GND\, F_BREADY => \GND\, F_RMW_AXI
         => \GND\, F_RREADY => \GND\, F_WDATA_HWDATA01(63) => 
        \VCC\, F_WDATA_HWDATA01(62) => \VCC\, 
        F_WDATA_HWDATA01(61) => \VCC\, F_WDATA_HWDATA01(60) => 
        \VCC\, F_WDATA_HWDATA01(59) => \VCC\, 
        F_WDATA_HWDATA01(58) => \VCC\, F_WDATA_HWDATA01(57) => 
        \VCC\, F_WDATA_HWDATA01(56) => \VCC\, 
        F_WDATA_HWDATA01(55) => \VCC\, F_WDATA_HWDATA01(54) => 
        \VCC\, F_WDATA_HWDATA01(53) => \VCC\, 
        F_WDATA_HWDATA01(52) => \VCC\, F_WDATA_HWDATA01(51) => 
        \VCC\, F_WDATA_HWDATA01(50) => \VCC\, 
        F_WDATA_HWDATA01(49) => \VCC\, F_WDATA_HWDATA01(48) => 
        \VCC\, F_WDATA_HWDATA01(47) => \VCC\, 
        F_WDATA_HWDATA01(46) => \VCC\, F_WDATA_HWDATA01(45) => 
        \VCC\, F_WDATA_HWDATA01(44) => \VCC\, 
        F_WDATA_HWDATA01(43) => \VCC\, F_WDATA_HWDATA01(42) => 
        \VCC\, F_WDATA_HWDATA01(41) => \VCC\, 
        F_WDATA_HWDATA01(40) => \VCC\, F_WDATA_HWDATA01(39) => 
        \VCC\, F_WDATA_HWDATA01(38) => \VCC\, 
        F_WDATA_HWDATA01(37) => \VCC\, F_WDATA_HWDATA01(36) => 
        \VCC\, F_WDATA_HWDATA01(35) => \VCC\, 
        F_WDATA_HWDATA01(34) => \VCC\, F_WDATA_HWDATA01(33) => 
        \VCC\, F_WDATA_HWDATA01(32) => \VCC\, 
        F_WDATA_HWDATA01(31) => \VCC\, F_WDATA_HWDATA01(30) => 
        \VCC\, F_WDATA_HWDATA01(29) => \VCC\, 
        F_WDATA_HWDATA01(28) => \VCC\, F_WDATA_HWDATA01(27) => 
        \VCC\, F_WDATA_HWDATA01(26) => \VCC\, 
        F_WDATA_HWDATA01(25) => \VCC\, F_WDATA_HWDATA01(24) => 
        \VCC\, F_WDATA_HWDATA01(23) => \VCC\, 
        F_WDATA_HWDATA01(22) => \VCC\, F_WDATA_HWDATA01(21) => 
        \VCC\, F_WDATA_HWDATA01(20) => \VCC\, 
        F_WDATA_HWDATA01(19) => \VCC\, F_WDATA_HWDATA01(18) => 
        \VCC\, F_WDATA_HWDATA01(17) => \VCC\, 
        F_WDATA_HWDATA01(16) => \VCC\, F_WDATA_HWDATA01(15) => 
        \VCC\, F_WDATA_HWDATA01(14) => \VCC\, 
        F_WDATA_HWDATA01(13) => \VCC\, F_WDATA_HWDATA01(12) => 
        \VCC\, F_WDATA_HWDATA01(11) => \VCC\, 
        F_WDATA_HWDATA01(10) => \VCC\, F_WDATA_HWDATA01(9) => 
        \VCC\, F_WDATA_HWDATA01(8) => \VCC\, F_WDATA_HWDATA01(7)
         => \VCC\, F_WDATA_HWDATA01(6) => \VCC\, 
        F_WDATA_HWDATA01(5) => \VCC\, F_WDATA_HWDATA01(4) => 
        \VCC\, F_WDATA_HWDATA01(3) => \VCC\, F_WDATA_HWDATA01(2)
         => \VCC\, F_WDATA_HWDATA01(1) => \VCC\, 
        F_WDATA_HWDATA01(0) => \VCC\, F_WID_HREADY01(3) => \GND\, 
        F_WID_HREADY01(2) => \GND\, F_WID_HREADY01(1) => \GND\, 
        F_WID_HREADY01(0) => \GND\, F_WLAST => \GND\, F_WSTRB(7)
         => \GND\, F_WSTRB(6) => \GND\, F_WSTRB(5) => \GND\, 
        F_WSTRB(4) => \GND\, F_WSTRB(3) => \GND\, F_WSTRB(2) => 
        \GND\, F_WSTRB(1) => \GND\, F_WSTRB(0) => \GND\, F_WVALID
         => \GND\, FPGA_MDDR_ARESET_N => \VCC\, 
        MDDR_FABRIC_PADDR(10) => \VCC\, MDDR_FABRIC_PADDR(9) => 
        \VCC\, MDDR_FABRIC_PADDR(8) => \VCC\, 
        MDDR_FABRIC_PADDR(7) => \VCC\, MDDR_FABRIC_PADDR(6) => 
        \VCC\, MDDR_FABRIC_PADDR(5) => \VCC\, 
        MDDR_FABRIC_PADDR(4) => \VCC\, MDDR_FABRIC_PADDR(3) => 
        \VCC\, MDDR_FABRIC_PADDR(2) => \VCC\, MDDR_FABRIC_PENABLE
         => \VCC\, MDDR_FABRIC_PSEL => \VCC\, 
        MDDR_FABRIC_PWDATA(15) => \VCC\, MDDR_FABRIC_PWDATA(14)
         => \VCC\, MDDR_FABRIC_PWDATA(13) => \VCC\, 
        MDDR_FABRIC_PWDATA(12) => \VCC\, MDDR_FABRIC_PWDATA(11)
         => \VCC\, MDDR_FABRIC_PWDATA(10) => \VCC\, 
        MDDR_FABRIC_PWDATA(9) => \VCC\, MDDR_FABRIC_PWDATA(8) => 
        \VCC\, MDDR_FABRIC_PWDATA(7) => \VCC\, 
        MDDR_FABRIC_PWDATA(6) => \VCC\, MDDR_FABRIC_PWDATA(5) => 
        \VCC\, MDDR_FABRIC_PWDATA(4) => \VCC\, 
        MDDR_FABRIC_PWDATA(3) => \VCC\, MDDR_FABRIC_PWDATA(2) => 
        \VCC\, MDDR_FABRIC_PWDATA(1) => \VCC\, 
        MDDR_FABRIC_PWDATA(0) => \VCC\, MDDR_FABRIC_PWRITE => 
        \VCC\, PRESET_N => \GND\, CAN_RXBUS_USBA_DATA1_MGPIO3A_IN
         => \GND\, CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => \GND\, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => \GND\, DM_IN(2) => 
        \GND\, DM_IN(1) => \GND\, DM_IN(0) => \GND\, 
        DRAM_DQ_IN(17) => \GND\, DRAM_DQ_IN(16) => \GND\, 
        DRAM_DQ_IN(15) => \GND\, DRAM_DQ_IN(14) => \GND\, 
        DRAM_DQ_IN(13) => \GND\, DRAM_DQ_IN(12) => \GND\, 
        DRAM_DQ_IN(11) => \GND\, DRAM_DQ_IN(10) => \GND\, 
        DRAM_DQ_IN(9) => \GND\, DRAM_DQ_IN(8) => \GND\, 
        DRAM_DQ_IN(7) => \GND\, DRAM_DQ_IN(6) => \GND\, 
        DRAM_DQ_IN(5) => \GND\, DRAM_DQ_IN(4) => \GND\, 
        DRAM_DQ_IN(3) => \GND\, DRAM_DQ_IN(2) => \GND\, 
        DRAM_DQ_IN(1) => \GND\, DRAM_DQ_IN(0) => \GND\, 
        DRAM_DQS_IN(2) => \GND\, DRAM_DQS_IN(1) => \GND\, 
        DRAM_DQS_IN(0) => \GND\, DRAM_FIFO_WE_IN(1) => \GND\, 
        DRAM_FIFO_WE_IN(0) => \GND\, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_IN => \GND\, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => \GND\, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => \GND\, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => \GND\, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => \GND\, 
        MMUART0_DCD_MGPIO22B_IN => \GND\, MMUART0_DSR_MGPIO20B_IN
         => \GND\, MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => \GND\, 
        MMUART0_RI_MGPIO21B_IN => \GND\, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => \GND\, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => MMUART_0_RXD_PAD_Y, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => \GND\, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => \GND\, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => MMUART_1_RXD_PAD_Y, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => \GND\, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => \GND\, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => \GND\, 
        RGMII_MDC_RMII_MDC_IN => \GND\, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => \GND\, 
        RGMII_RX_CLK_IN => \GND\, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => \GND\, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => \GND\, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => \GND\, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => \GND\, 
        RGMII_RXD3_USBB_DATA4_IN => \GND\, RGMII_TX_CLK_IN => 
        \GND\, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => \GND\, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => \GND\, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => \GND\, 
        RGMII_TXD2_USBB_DATA5_IN => \GND\, 
        RGMII_TXD3_USBB_DATA6_IN => \GND\, SPI0_SCK_USBA_XCLK_IN
         => \GND\, SPI0_SDI_USBA_DIR_MGPIO5A_IN => \GND\, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => \GND\, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => \GND\, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => \GND\, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => \GND\, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => \GND\, SPI1_SCK_IN => 
        \GND\, SPI1_SDI_MGPIO11A_IN => \GND\, 
        SPI1_SDO_MGPIO12A_IN => \GND\, SPI1_SS0_MGPIO13A_IN => 
        \GND\, SPI1_SS1_MGPIO14A_IN => \GND\, 
        SPI1_SS2_MGPIO15A_IN => \GND\, SPI1_SS3_MGPIO16A_IN => 
        \GND\, SPI1_SS4_MGPIO17A_IN => \GND\, 
        SPI1_SS5_MGPIO18A_IN => \GND\, SPI1_SS6_MGPIO23A_IN => 
        \GND\, SPI1_SS7_MGPIO24A_IN => \GND\, USBC_XCLK_IN => 
        \GND\, CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT, DRAM_ADDR(15) => 
        DRAM_ADDR(15), DRAM_ADDR(14) => DRAM_ADDR(14), 
        DRAM_ADDR(13) => DRAM_ADDR(13), DRAM_ADDR(12) => 
        DRAM_ADDR(12), DRAM_ADDR(11) => DRAM_ADDR(11), 
        DRAM_ADDR(10) => DRAM_ADDR(10), DRAM_ADDR(9) => 
        DRAM_ADDR(9), DRAM_ADDR(8) => DRAM_ADDR(8), DRAM_ADDR(7)
         => DRAM_ADDR(7), DRAM_ADDR(6) => DRAM_ADDR(6), 
        DRAM_ADDR(5) => DRAM_ADDR(5), DRAM_ADDR(4) => 
        DRAM_ADDR(4), DRAM_ADDR(3) => DRAM_ADDR(3), DRAM_ADDR(2)
         => DRAM_ADDR(2), DRAM_ADDR(1) => DRAM_ADDR(1), 
        DRAM_ADDR(0) => DRAM_ADDR(0), DRAM_BA(2) => DRAM_BA(2), 
        DRAM_BA(1) => DRAM_BA(1), DRAM_BA(0) => DRAM_BA(0), 
        DRAM_CASN => DRAM_CASN, DRAM_CKE => DRAM_CKE, DRAM_CLK
         => DRAM_CLK, DRAM_CSN => DRAM_CSN, DRAM_DM_RDQS_OUT(2)
         => DRAM_DM_RDQS_OUT(2), DRAM_DM_RDQS_OUT(1) => 
        DRAM_DM_RDQS_OUT(1), DRAM_DM_RDQS_OUT(0) => 
        DRAM_DM_RDQS_OUT(0), DRAM_DQ_OUT(17) => DRAM_DQ_OUT(17), 
        DRAM_DQ_OUT(16) => DRAM_DQ_OUT(16), DRAM_DQ_OUT(15) => 
        DRAM_DQ_OUT(15), DRAM_DQ_OUT(14) => DRAM_DQ_OUT(14), 
        DRAM_DQ_OUT(13) => DRAM_DQ_OUT(13), DRAM_DQ_OUT(12) => 
        DRAM_DQ_OUT(12), DRAM_DQ_OUT(11) => DRAM_DQ_OUT(11), 
        DRAM_DQ_OUT(10) => DRAM_DQ_OUT(10), DRAM_DQ_OUT(9) => 
        DRAM_DQ_OUT(9), DRAM_DQ_OUT(8) => DRAM_DQ_OUT(8), 
        DRAM_DQ_OUT(7) => DRAM_DQ_OUT(7), DRAM_DQ_OUT(6) => 
        DRAM_DQ_OUT(6), DRAM_DQ_OUT(5) => DRAM_DQ_OUT(5), 
        DRAM_DQ_OUT(4) => DRAM_DQ_OUT(4), DRAM_DQ_OUT(3) => 
        DRAM_DQ_OUT(3), DRAM_DQ_OUT(2) => DRAM_DQ_OUT(2), 
        DRAM_DQ_OUT(1) => DRAM_DQ_OUT(1), DRAM_DQ_OUT(0) => 
        DRAM_DQ_OUT(0), DRAM_DQS_OUT(2) => DRAM_DQS_OUT(2), 
        DRAM_DQS_OUT(1) => DRAM_DQS_OUT(1), DRAM_DQS_OUT(0) => 
        DRAM_DQS_OUT(0), DRAM_FIFO_WE_OUT(1) => 
        DRAM_FIFO_WE_OUT(1), DRAM_FIFO_WE_OUT(0) => 
        DRAM_FIFO_WE_OUT(0), DRAM_ODT => DRAM_ODT, DRAM_RASN => 
        DRAM_RASN, DRAM_RSTN => DRAM_RSTN, DRAM_WEN => DRAM_WEN, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OUT => 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OUT, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OUT, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT => 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT, 
        MMUART0_DCD_MGPIO22B_OUT => MMUART0_DCD_MGPIO22B_OUT, 
        MMUART0_DSR_MGPIO20B_OUT => MMUART0_DSR_MGPIO20B_OUT, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT, 
        MMUART0_RI_MGPIO21B_OUT => MMUART0_RI_MGPIO21B_OUT, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT, 
        RGMII_MDC_RMII_MDC_OUT => RGMII_MDC_RMII_MDC_OUT, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT, RGMII_RX_CLK_OUT => 
        RGMII_RX_CLK_OUT, RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT
         => RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT, 
        RGMII_RXD3_USBB_DATA4_OUT => RGMII_RXD3_USBB_DATA4_OUT, 
        RGMII_TX_CLK_OUT => RGMII_TX_CLK_OUT, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT, 
        RGMII_TXD2_USBB_DATA5_OUT => RGMII_TXD2_USBB_DATA5_OUT, 
        RGMII_TXD3_USBB_DATA6_OUT => RGMII_TXD3_USBB_DATA6_OUT, 
        SPI0_SCK_USBA_XCLK_OUT => SPI0_SCK_USBA_XCLK_OUT, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT => 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT, SPI1_SCK_OUT => 
        SPI1_SCK_OUT, SPI1_SDI_MGPIO11A_OUT => 
        SPI1_SDI_MGPIO11A_OUT, SPI1_SDO_MGPIO12A_OUT => 
        SPI1_SDO_MGPIO12A_OUT, SPI1_SS0_MGPIO13A_OUT => 
        SPI1_SS0_MGPIO13A_OUT, SPI1_SS1_MGPIO14A_OUT => 
        SPI1_SS1_MGPIO14A_OUT, SPI1_SS2_MGPIO15A_OUT => 
        SPI1_SS2_MGPIO15A_OUT, SPI1_SS3_MGPIO16A_OUT => 
        SPI1_SS3_MGPIO16A_OUT, SPI1_SS4_MGPIO17A_OUT => 
        SPI1_SS4_MGPIO17A_OUT, SPI1_SS5_MGPIO18A_OUT => 
        SPI1_SS5_MGPIO18A_OUT, SPI1_SS6_MGPIO23A_OUT => 
        SPI1_SS6_MGPIO23A_OUT, SPI1_SS7_MGPIO24A_OUT => 
        SPI1_SS7_MGPIO24A_OUT, USBC_XCLK_OUT => USBC_XCLK_OUT, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE, DM_OE(2) => DM_OE(2), 
        DM_OE(1) => DM_OE(1), DM_OE(0) => DM_OE(0), 
        DRAM_DQ_OE(17) => DRAM_DQ_OE(17), DRAM_DQ_OE(16) => 
        DRAM_DQ_OE(16), DRAM_DQ_OE(15) => DRAM_DQ_OE(15), 
        DRAM_DQ_OE(14) => DRAM_DQ_OE(14), DRAM_DQ_OE(13) => 
        DRAM_DQ_OE(13), DRAM_DQ_OE(12) => DRAM_DQ_OE(12), 
        DRAM_DQ_OE(11) => DRAM_DQ_OE(11), DRAM_DQ_OE(10) => 
        DRAM_DQ_OE(10), DRAM_DQ_OE(9) => DRAM_DQ_OE(9), 
        DRAM_DQ_OE(8) => DRAM_DQ_OE(8), DRAM_DQ_OE(7) => 
        DRAM_DQ_OE(7), DRAM_DQ_OE(6) => DRAM_DQ_OE(6), 
        DRAM_DQ_OE(5) => DRAM_DQ_OE(5), DRAM_DQ_OE(4) => 
        DRAM_DQ_OE(4), DRAM_DQ_OE(3) => DRAM_DQ_OE(3), 
        DRAM_DQ_OE(2) => DRAM_DQ_OE(2), DRAM_DQ_OE(1) => 
        DRAM_DQ_OE(1), DRAM_DQ_OE(0) => DRAM_DQ_OE(0), 
        DRAM_DQS_OE(2) => DRAM_DQS_OE(2), DRAM_DQS_OE(1) => 
        DRAM_DQS_OE(1), DRAM_DQS_OE(0) => DRAM_DQS_OE(0), 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE => 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE, 
        MMUART0_DCD_MGPIO22B_OE => MMUART0_DCD_MGPIO22B_OE, 
        MMUART0_DSR_MGPIO20B_OE => MMUART0_DSR_MGPIO20B_OE, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OE, 
        MMUART0_RI_MGPIO21B_OE => MMUART0_RI_MGPIO21B_OE, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE, 
        RGMII_MDC_RMII_MDC_OE => RGMII_MDC_RMII_MDC_OE, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE, RGMII_RX_CLK_OE => 
        RGMII_RX_CLK_OE, RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE
         => RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE, 
        RGMII_RXD3_USBB_DATA4_OE => RGMII_RXD3_USBB_DATA4_OE, 
        RGMII_TX_CLK_OE => RGMII_TX_CLK_OE, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE, 
        RGMII_TXD2_USBB_DATA5_OE => RGMII_TXD2_USBB_DATA5_OE, 
        RGMII_TXD3_USBB_DATA6_OE => RGMII_TXD3_USBB_DATA6_OE, 
        SPI0_SCK_USBA_XCLK_OE => SPI0_SCK_USBA_XCLK_OE, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OE => 
        SPI0_SDI_USBA_DIR_MGPIO5A_OE, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => 
        SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE, SPI1_SCK_OE => 
        SPI1_SCK_OE, SPI1_SDI_MGPIO11A_OE => SPI1_SDI_MGPIO11A_OE, 
        SPI1_SDO_MGPIO12A_OE => SPI1_SDO_MGPIO12A_OE, 
        SPI1_SS0_MGPIO13A_OE => SPI1_SS0_MGPIO13A_OE, 
        SPI1_SS1_MGPIO14A_OE => SPI1_SS1_MGPIO14A_OE, 
        SPI1_SS2_MGPIO15A_OE => SPI1_SS2_MGPIO15A_OE, 
        SPI1_SS3_MGPIO16A_OE => SPI1_SS3_MGPIO16A_OE, 
        SPI1_SS4_MGPIO17A_OE => SPI1_SS4_MGPIO17A_OE, 
        SPI1_SS5_MGPIO18A_OE => SPI1_SS5_MGPIO18A_OE, 
        SPI1_SS6_MGPIO23A_OE => SPI1_SS6_MGPIO23A_OE, 
        SPI1_SS7_MGPIO24A_OE => SPI1_SS7_MGPIO24A_OE, 
        USBC_XCLK_OE => USBC_XCLK_OE);
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    MMUART_1_TXD_PAD : TRIBUFF
      generic map(IOSTD => "")

      port map(D => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, PAD
         => TM_TX);
    
    MMUART_1_RXD_PAD : INBUF
      generic map(IOSTD => "")

      port map(PAD => TM_RX, Y => MMUART_1_RXD_PAD_Y);
    
    MMUART_0_TXD_PAD : TRIBUFF
      generic map(IOSTD => "")

      port map(D => 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, E => 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, PAD => 
        DAPI_TX);
    
    GND_Z : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sb_sb_FABOSC_0_OSC is

    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );

end sb_sb_FABOSC_0_OSC;

architecture DEF_ARCH of sb_sb_FABOSC_0_OSC is 

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \GND\, \VCC\ : std_logic;

begin 


    I_RCOSC_25_50MHZ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.000000)

      port map(CLKOUT => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    GND_Z : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAPB3_MUXPTOB3 is

    port( sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : out   std_logic_vector(31 downto 0);
          sb_sb_0_Memory_PRDATA                   : in    std_logic_vector(31 downto 0);
          sb_sb_0_STAMP_PRDATA                    : in    std_logic_vector(31 downto 0);
          STAMP_PADDRS                            : in    std_logic_vector(14 downto 12);
          iPSELS_raw_1_0                          : in    std_logic;
          PRDATA_N_5_i                            : out   std_logic;
          sb_sb_0_Memory_PREADY                   : in    std_logic;
          sb_sb_0_STAMP_PREADY                    : in    std_logic;
          PREADY_N_7                              : out   std_logic;
          sb_sb_0_Memory_PSELx                    : in    std_logic
        );

end COREAPB3_MUXPTOB3;

architecture DEF_ARCH of COREAPB3_MUXPTOB3 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal PSELSBUS_Z : std_logic_vector(2 downto 0);
    signal PSELSBUS : std_logic_vector(1 to 1);
    signal PRDATA_0_iv_1 : std_logic_vector(0 to 0);
    signal PREADY_m4_i_sx_Z, iprdata46_Z, PRDATA_N_7, \GND\, 
        \VCC\ : std_logic;

begin 


    \PRDATA_0_iv[12]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(12), B => 
        sb_sb_0_Memory_PRDATA(12), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12));
    
    \PRDATA_0_iv[19]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(19), B => 
        sb_sb_0_Memory_PRDATA(19), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19));
    
    iPRDATA_0_sqmuxa : CFG4
      generic map(INIT => x"0002")

      port map(A => sb_sb_0_Memory_PSELx, B => PSELSBUS_Z(0), C
         => PSELSBUS_Z(2), D => PSELSBUS(1), Y => 
        PRDATA_0_iv_1(0));
    
    \PSELSBUS[2]\ : CFG4
      generic map(INIT => x"20A0")

      port map(A => STAMP_PADDRS(14), B => STAMP_PADDRS(13), C
         => iPSELS_raw_1_0, D => STAMP_PADDRS(12), Y => 
        PSELSBUS_Z(2));
    
    \PRDATA_0_iv[18]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(18), B => 
        sb_sb_0_Memory_PRDATA(18), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18));
    
    \PRDATA_0_iv[16]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(16), B => 
        sb_sb_0_Memory_PRDATA(16), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16));
    
    \PRDATA_0_iv[11]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(11), B => 
        sb_sb_0_Memory_PRDATA(11), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11));
    
    \PRDATA_0_iv[10]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(10), B => 
        sb_sb_0_Memory_PRDATA(10), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10));
    
    \PRDATA_0_iv[0]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(0), B => 
        sb_sb_0_Memory_PRDATA(0), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(0));
    
    \PSELSBUS_1[1]\ : CFG4
      generic map(INIT => x"40C0")

      port map(A => STAMP_PADDRS(14), B => STAMP_PADDRS(13), C
         => iPSELS_raw_1_0, D => STAMP_PADDRS(12), Y => 
        PSELSBUS(1));
    
    \PRDATA_0_iv[14]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(14), B => 
        sb_sb_0_Memory_PRDATA(14), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14));
    
    \PRDATA_0_iv[2]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(2), B => 
        sb_sb_0_Memory_PRDATA(2), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(2));
    
    \PRDATA_0_iv[9]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(9), B => 
        sb_sb_0_Memory_PRDATA(9), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9));
    
    \PRDATA_0_iv[5]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(5), B => 
        sb_sb_0_Memory_PRDATA(5), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(5));
    
    \PRDATA_0_iv[22]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(22), B => 
        sb_sb_0_Memory_PRDATA(22), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22));
    
    \PRDATA_0_iv[13]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(13), B => 
        sb_sb_0_Memory_PRDATA(13), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13));
    
    \PRDATA_0_iv[29]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(29), B => 
        sb_sb_0_Memory_PRDATA(29), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29));
    
    \PRDATA_0_iv[15]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(15), B => 
        sb_sb_0_Memory_PRDATA(15), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15));
    
    \PRDATA_0_iv[17]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(17), B => 
        sb_sb_0_Memory_PRDATA(17), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17));
    
    \PRDATA_0_iv[4]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(4), B => 
        sb_sb_0_Memory_PRDATA(4), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(4));
    
    PRDATA_m4_0_m3 : CFG4
      generic map(INIT => x"AAC0")

      port map(A => sb_sb_0_STAMP_PRDATA(3), B => 
        sb_sb_0_Memory_PRDATA(3), C => sb_sb_0_Memory_PSELx, D
         => PSELSBUS_Z(0), Y => PRDATA_N_7);
    
    iprdata46 : CFG3
      generic map(INIT => x"10")

      port map(A => PSELSBUS_Z(2), B => PSELSBUS(1), C => 
        PSELSBUS_Z(0), Y => iprdata46_Z);
    
    \PRDATA_0_iv[28]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(28), B => 
        sb_sb_0_Memory_PRDATA(28), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28));
    
    \PRDATA_0_iv[26]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(26), B => 
        sb_sb_0_Memory_PRDATA(26), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26));
    
    \PRDATA_0_iv[1]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(1), B => 
        sb_sb_0_Memory_PRDATA(1), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(1));
    
    \PRDATA_0_iv[21]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(21), B => 
        sb_sb_0_Memory_PRDATA(21), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21));
    
    \PRDATA_0_iv[20]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(20), B => 
        sb_sb_0_Memory_PRDATA(20), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20));
    
    \PRDATA_0_iv[8]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(8), B => 
        sb_sb_0_Memory_PRDATA(8), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8));
    
    \PRDATA_0_iv[6]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(6), B => 
        sb_sb_0_Memory_PRDATA(6), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(6));
    
    \PRDATA_0_iv[24]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(24), B => 
        sb_sb_0_Memory_PRDATA(24), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24));
    
    \PRDATA_0_iv[7]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(7), B => 
        sb_sb_0_Memory_PRDATA(7), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(7));
    
    PREADY_m4_i_sx : CFG4
      generic map(INIT => x"FAFC")

      port map(A => sb_sb_0_STAMP_PREADY, B => 
        sb_sb_0_Memory_PREADY, C => PSELSBUS(1), D => 
        PSELSBUS_Z(0), Y => PREADY_m4_i_sx_Z);
    
    GND_Z : GND
      port map(Y => \GND\);
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    \PSELSBUS[0]\ : CFG4
      generic map(INIT => x"7000")

      port map(A => STAMP_PADDRS(14), B => STAMP_PADDRS(13), C
         => iPSELS_raw_1_0, D => STAMP_PADDRS(12), Y => 
        PSELSBUS_Z(0));
    
    \PRDATA_0_iv[31]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(31), B => 
        sb_sb_0_Memory_PRDATA(31), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31));
    
    \PRDATA_0_iv[30]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(30), B => 
        sb_sb_0_Memory_PRDATA(30), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30));
    
    \PRDATA_0_iv[23]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(23), B => 
        sb_sb_0_Memory_PRDATA(23), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23));
    
    \PRDATA_0_iv[25]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(25), B => 
        sb_sb_0_Memory_PRDATA(25), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25));
    
    \PRDATA_0_iv[27]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => sb_sb_0_STAMP_PRDATA(27), B => 
        sb_sb_0_Memory_PRDATA(27), C => iprdata46_Z, D => 
        PRDATA_0_iv_1(0), Y => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27));
    
    PREADY_m4_i : CFG4
      generic map(INIT => x"FCFD")

      port map(A => sb_sb_0_Memory_PSELx, B => PSELSBUS_Z(2), C
         => PREADY_m4_i_sx_Z, D => PSELSBUS_Z(0), Y => PREADY_N_7);
    
    PRDATA_m4_0_m3_RNI8EAL : CFG3
      generic map(INIT => x"10")

      port map(A => PSELSBUS_Z(2), B => PSELSBUS(1), C => 
        PRDATA_N_7, Y => PRDATA_N_5_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAPB3 is

    port( sb_sb_0_STAMP_PRDATA                    : in    std_logic_vector(31 downto 0);
          sb_sb_0_Memory_PRDATA                   : in    std_logic_vector(31 downto 0);
          sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : out   std_logic_vector(31 downto 0);
          STAMP_PADDRS                            : in    std_logic_vector(15 downto 12);
          PREADY_N_7                              : out   std_logic;
          sb_sb_0_STAMP_PREADY                    : in    std_logic;
          sb_sb_0_Memory_PREADY                   : in    std_logic;
          PRDATA_N_5_i                            : out   std_logic;
          sb_sb_0_STAMP_PSELx                     : out   std_logic;
          sb_sb_0_Memory_PSELx                    : out   std_logic;
          sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx  : in    std_logic
        );

end CoreAPB3;

architecture DEF_ARCH of CoreAPB3 is 

  component COREAPB3_MUXPTOB3
    port( sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : out   std_logic_vector(31 downto 0);
          sb_sb_0_Memory_PRDATA                   : in    std_logic_vector(31 downto 0) := (others => 'U');
          sb_sb_0_STAMP_PRDATA                    : in    std_logic_vector(31 downto 0) := (others => 'U');
          STAMP_PADDRS                            : in    std_logic_vector(14 downto 12) := (others => 'U');
          iPSELS_raw_1_0                          : in    std_logic := 'U';
          PRDATA_N_5_i                            : out   std_logic;
          sb_sb_0_Memory_PREADY                   : in    std_logic := 'U';
          sb_sb_0_STAMP_PREADY                    : in    std_logic := 'U';
          PREADY_N_7                              : out   std_logic;
          sb_sb_0_Memory_PSELx                    : in    std_logic := 'U'
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \sb_sb_0_Memory_PSELx\ : std_logic;
    signal iPSELS_raw_1 : std_logic_vector(0 to 0);
    signal N_2041, \GND\, \VCC\ : std_logic;

    for all : COREAPB3_MUXPTOB3
	Use entity work.COREAPB3_MUXPTOB3(DEF_ARCH);
begin 

    sb_sb_0_Memory_PSELx <= \sb_sb_0_Memory_PSELx\;

    u_mux_p_to_b3 : COREAPB3_MUXPTOB3
      port map(sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(7) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(7), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(6) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(6), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(5) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(5), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(4) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(4), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(3) => N_2041, 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(2) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(2), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(1) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(1), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(0) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(0), 
        sb_sb_0_Memory_PRDATA(31) => sb_sb_0_Memory_PRDATA(31), 
        sb_sb_0_Memory_PRDATA(30) => sb_sb_0_Memory_PRDATA(30), 
        sb_sb_0_Memory_PRDATA(29) => sb_sb_0_Memory_PRDATA(29), 
        sb_sb_0_Memory_PRDATA(28) => sb_sb_0_Memory_PRDATA(28), 
        sb_sb_0_Memory_PRDATA(27) => sb_sb_0_Memory_PRDATA(27), 
        sb_sb_0_Memory_PRDATA(26) => sb_sb_0_Memory_PRDATA(26), 
        sb_sb_0_Memory_PRDATA(25) => sb_sb_0_Memory_PRDATA(25), 
        sb_sb_0_Memory_PRDATA(24) => sb_sb_0_Memory_PRDATA(24), 
        sb_sb_0_Memory_PRDATA(23) => sb_sb_0_Memory_PRDATA(23), 
        sb_sb_0_Memory_PRDATA(22) => sb_sb_0_Memory_PRDATA(22), 
        sb_sb_0_Memory_PRDATA(21) => sb_sb_0_Memory_PRDATA(21), 
        sb_sb_0_Memory_PRDATA(20) => sb_sb_0_Memory_PRDATA(20), 
        sb_sb_0_Memory_PRDATA(19) => sb_sb_0_Memory_PRDATA(19), 
        sb_sb_0_Memory_PRDATA(18) => sb_sb_0_Memory_PRDATA(18), 
        sb_sb_0_Memory_PRDATA(17) => sb_sb_0_Memory_PRDATA(17), 
        sb_sb_0_Memory_PRDATA(16) => sb_sb_0_Memory_PRDATA(16), 
        sb_sb_0_Memory_PRDATA(15) => sb_sb_0_Memory_PRDATA(15), 
        sb_sb_0_Memory_PRDATA(14) => sb_sb_0_Memory_PRDATA(14), 
        sb_sb_0_Memory_PRDATA(13) => sb_sb_0_Memory_PRDATA(13), 
        sb_sb_0_Memory_PRDATA(12) => sb_sb_0_Memory_PRDATA(12), 
        sb_sb_0_Memory_PRDATA(11) => sb_sb_0_Memory_PRDATA(11), 
        sb_sb_0_Memory_PRDATA(10) => sb_sb_0_Memory_PRDATA(10), 
        sb_sb_0_Memory_PRDATA(9) => sb_sb_0_Memory_PRDATA(9), 
        sb_sb_0_Memory_PRDATA(8) => sb_sb_0_Memory_PRDATA(8), 
        sb_sb_0_Memory_PRDATA(7) => sb_sb_0_Memory_PRDATA(7), 
        sb_sb_0_Memory_PRDATA(6) => sb_sb_0_Memory_PRDATA(6), 
        sb_sb_0_Memory_PRDATA(5) => sb_sb_0_Memory_PRDATA(5), 
        sb_sb_0_Memory_PRDATA(4) => sb_sb_0_Memory_PRDATA(4), 
        sb_sb_0_Memory_PRDATA(3) => sb_sb_0_Memory_PRDATA(3), 
        sb_sb_0_Memory_PRDATA(2) => sb_sb_0_Memory_PRDATA(2), 
        sb_sb_0_Memory_PRDATA(1) => sb_sb_0_Memory_PRDATA(1), 
        sb_sb_0_Memory_PRDATA(0) => sb_sb_0_Memory_PRDATA(0), 
        sb_sb_0_STAMP_PRDATA(31) => sb_sb_0_STAMP_PRDATA(31), 
        sb_sb_0_STAMP_PRDATA(30) => sb_sb_0_STAMP_PRDATA(30), 
        sb_sb_0_STAMP_PRDATA(29) => sb_sb_0_STAMP_PRDATA(29), 
        sb_sb_0_STAMP_PRDATA(28) => sb_sb_0_STAMP_PRDATA(28), 
        sb_sb_0_STAMP_PRDATA(27) => sb_sb_0_STAMP_PRDATA(27), 
        sb_sb_0_STAMP_PRDATA(26) => sb_sb_0_STAMP_PRDATA(26), 
        sb_sb_0_STAMP_PRDATA(25) => sb_sb_0_STAMP_PRDATA(25), 
        sb_sb_0_STAMP_PRDATA(24) => sb_sb_0_STAMP_PRDATA(24), 
        sb_sb_0_STAMP_PRDATA(23) => sb_sb_0_STAMP_PRDATA(23), 
        sb_sb_0_STAMP_PRDATA(22) => sb_sb_0_STAMP_PRDATA(22), 
        sb_sb_0_STAMP_PRDATA(21) => sb_sb_0_STAMP_PRDATA(21), 
        sb_sb_0_STAMP_PRDATA(20) => sb_sb_0_STAMP_PRDATA(20), 
        sb_sb_0_STAMP_PRDATA(19) => sb_sb_0_STAMP_PRDATA(19), 
        sb_sb_0_STAMP_PRDATA(18) => sb_sb_0_STAMP_PRDATA(18), 
        sb_sb_0_STAMP_PRDATA(17) => sb_sb_0_STAMP_PRDATA(17), 
        sb_sb_0_STAMP_PRDATA(16) => sb_sb_0_STAMP_PRDATA(16), 
        sb_sb_0_STAMP_PRDATA(15) => sb_sb_0_STAMP_PRDATA(15), 
        sb_sb_0_STAMP_PRDATA(14) => sb_sb_0_STAMP_PRDATA(14), 
        sb_sb_0_STAMP_PRDATA(13) => sb_sb_0_STAMP_PRDATA(13), 
        sb_sb_0_STAMP_PRDATA(12) => sb_sb_0_STAMP_PRDATA(12), 
        sb_sb_0_STAMP_PRDATA(11) => sb_sb_0_STAMP_PRDATA(11), 
        sb_sb_0_STAMP_PRDATA(10) => sb_sb_0_STAMP_PRDATA(10), 
        sb_sb_0_STAMP_PRDATA(9) => sb_sb_0_STAMP_PRDATA(9), 
        sb_sb_0_STAMP_PRDATA(8) => sb_sb_0_STAMP_PRDATA(8), 
        sb_sb_0_STAMP_PRDATA(7) => sb_sb_0_STAMP_PRDATA(7), 
        sb_sb_0_STAMP_PRDATA(6) => sb_sb_0_STAMP_PRDATA(6), 
        sb_sb_0_STAMP_PRDATA(5) => sb_sb_0_STAMP_PRDATA(5), 
        sb_sb_0_STAMP_PRDATA(4) => sb_sb_0_STAMP_PRDATA(4), 
        sb_sb_0_STAMP_PRDATA(3) => sb_sb_0_STAMP_PRDATA(3), 
        sb_sb_0_STAMP_PRDATA(2) => sb_sb_0_STAMP_PRDATA(2), 
        sb_sb_0_STAMP_PRDATA(1) => sb_sb_0_STAMP_PRDATA(1), 
        sb_sb_0_STAMP_PRDATA(0) => sb_sb_0_STAMP_PRDATA(0), 
        STAMP_PADDRS(14) => STAMP_PADDRS(14), STAMP_PADDRS(13)
         => STAMP_PADDRS(13), STAMP_PADDRS(12) => 
        STAMP_PADDRS(12), iPSELS_raw_1_0 => iPSELS_raw_1(0), 
        PRDATA_N_5_i => PRDATA_N_5_i, sb_sb_0_Memory_PREADY => 
        sb_sb_0_Memory_PREADY, sb_sb_0_STAMP_PREADY => 
        sb_sb_0_STAMP_PREADY, PREADY_N_7 => PREADY_N_7, 
        sb_sb_0_Memory_PSELx => \sb_sb_0_Memory_PSELx\);
    
    \iPSELS_raw_1_0[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => STAMP_PADDRS(15), B => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, Y => 
        iPSELS_raw_1(0));
    
    \iPSELS_raw[1]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => STAMP_PADDRS(14), B => STAMP_PADDRS(13), C
         => iPSELS_raw_1(0), D => STAMP_PADDRS(12), Y => 
        sb_sb_0_STAMP_PSELx);
    
    \iPSELS_raw[0]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => STAMP_PADDRS(14), B => STAMP_PADDRS(13), C
         => iPSELS_raw_1(0), D => STAMP_PADDRS(12), Y => 
        \sb_sb_0_Memory_PSELx\);
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    GND_Z : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sb_sb_CCC_0_FCCC is

    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic;
          FIC_0_LOCK                                         : out   std_logic;
          adc_clk_c                                          : out   std_logic;
          sb_sb_0_FIC_0_CLK                                  : out   std_logic
        );

end sb_sb_CCC_0_FCCC;

architecture DEF_ARCH of sb_sb_CCC_0_FCCC is 

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal PRDATA : std_logic_vector(7 downto 0);
    signal GL0_net, GL1_net, Y0, Y1, Y2, Y3, BUSY, \VCC\, \GND\, 
        GL2, GL3 : std_logic;

begin 


    GL1_INST : CLKINT
      port map(A => GL1_net, Y => adc_clk_c);
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => sb_sb_0_FIC_0_CLK);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FB8000044174000F18C6309C231839DEC0407A04C02501",
         VCOFREQUENCY => 950.000000)

      port map(Y0 => Y0, Y1 => Y1, Y2 => Y2, Y3 => Y3, PRDATA(7)
         => PRDATA(7), PRDATA(6) => PRDATA(6), PRDATA(5) => 
        PRDATA(5), PRDATA(4) => PRDATA(4), PRDATA(3) => PRDATA(3), 
        PRDATA(2) => PRDATA(2), PRDATA(1) => PRDATA(1), PRDATA(0)
         => PRDATA(0), LOCK => FIC_0_LOCK, BUSY => BUSY, CLK0 => 
        \VCC\, CLK1 => \VCC\, CLK2 => \VCC\, CLK3 => \VCC\, 
        NGMUX0_SEL => \GND\, NGMUX1_SEL => \GND\, NGMUX2_SEL => 
        \GND\, NGMUX3_SEL => \GND\, NGMUX0_HOLD_N => \VCC\, 
        NGMUX1_HOLD_N => \VCC\, NGMUX2_HOLD_N => \VCC\, 
        NGMUX3_HOLD_N => \VCC\, NGMUX0_ARST_N => \VCC\, 
        NGMUX1_ARST_N => \VCC\, NGMUX2_ARST_N => \VCC\, 
        NGMUX3_ARST_N => \VCC\, PLL_BYPASS_N => \VCC\, PLL_ARST_N
         => \VCC\, PLL_POWERDOWN_N => \VCC\, GPD0_ARST_N => \VCC\, 
        GPD1_ARST_N => \VCC\, GPD2_ARST_N => \VCC\, GPD3_ARST_N
         => \VCC\, PRESET_N => \GND\, PCLK => \VCC\, PSEL => 
        \VCC\, PENABLE => \VCC\, PWRITE => \VCC\, PADDR(7) => 
        \VCC\, PADDR(6) => \VCC\, PADDR(5) => \VCC\, PADDR(4) => 
        \VCC\, PADDR(3) => \VCC\, PADDR(2) => \VCC\, PWDATA(7)
         => \VCC\, PWDATA(6) => \VCC\, PWDATA(5) => \VCC\, 
        PWDATA(4) => \VCC\, PWDATA(3) => \VCC\, PWDATA(2) => 
        \VCC\, PWDATA(1) => \VCC\, PWDATA(0) => \VCC\, CLK0_PAD
         => \GND\, CLK1_PAD => \GND\, CLK2_PAD => \GND\, CLK3_PAD
         => \GND\, GL0 => GL0_net, GL1 => GL1_net, GL2 => GL2, 
        GL3 => GL3, RCOSC_25_50MHZ => 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        RCOSC_1MHZ => \GND\, XTLOSC => \GND\);
    
    GND_Z : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sb_sb is

    port( sb_sb_0_STAMP_PADDR      : out   std_logic_vector(11 downto 0);
          sb_sb_0_STAMP_PWDATA     : out   std_logic_vector(31 downto 0);
          dataReady_0              : in    std_logic;
          sb_sb_0_Memory_PRDATA    : in    std_logic_vector(31 downto 0);
          sb_sb_0_STAMP_PRDATA     : in    std_logic_vector(31 downto 0);
          TM_TX                    : out   std_logic;
          TM_RX                    : in    std_logic;
          DAPI_TX                  : out   std_logic;
          DAPI_RX                  : in    std_logic;
          sb_sb_0_GPIO_3_M2F       : out   std_logic;
          sb_sb_0_GPIO_4_M2F       : out   std_logic;
          sb_sb_0_STAMP_PENABLE    : out   std_logic;
          sb_sb_0_STAMP_PWRITE     : out   std_logic;
          LED_HEARTBEAT_c          : out   std_logic;
          LED_RECORDING_c          : out   std_logic;
          GPIO_6_M2F_c             : out   std_logic;
          RXSM_LO_c                : in    std_logic;
          RXSM_SOE_c               : in    std_logic;
          RXSM_SODS_c              : in    std_logic;
          sb_sb_0_Memory_PSELx     : out   std_logic;
          sb_sb_0_STAMP_PSELx      : out   std_logic;
          sb_sb_0_Memory_PREADY    : in    std_logic;
          sb_sb_0_STAMP_PREADY     : in    std_logic;
          sb_sb_0_FIC_0_CLK        : out   std_logic;
          adc_clk_c                : out   std_logic;
          DEVRST_N                 : in    std_logic;
          sb_sb_0_POWER_ON_RESET_N : out   std_logic
        );

end sb_sb;

architecture DEF_ARCH of sb_sb is 

  component sb_sb_MSS
    port( sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : in    std_logic_vector(31 downto 0) := (others => 'U');
          dataReady_0                             : in    std_logic := 'U';
          sb_sb_0_STAMP_PWDATA                    : out   std_logic_vector(31 downto 0);
          STAMP_PADDRS                            : out   std_logic_vector(15 downto 12);
          sb_sb_0_STAMP_PADDR                     : out   std_logic_vector(11 downto 0);
          sb_sb_0_FIC_0_CLK                       : in    std_logic := 'U';
          RXSM_SODS_c                             : in    std_logic := 'U';
          RXSM_SOE_c                              : in    std_logic := 'U';
          RXSM_LO_c                               : in    std_logic := 'U';
          FIC_0_LOCK                              : in    std_logic := 'U';
          PREADY_N_7                              : in    std_logic := 'U';
          PRDATA_N_5_i                            : in    std_logic := 'U';
          GPIO_6_M2F_c                            : out   std_logic;
          LED_RECORDING_c                         : out   std_logic;
          LED_HEARTBEAT_c                         : out   std_logic;
          sb_sb_0_STAMP_PWRITE                    : out   std_logic;
          sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx  : out   std_logic;
          sb_sb_0_STAMP_PENABLE                   : out   std_logic;
          sb_sb_0_GPIO_4_M2F                      : out   std_logic;
          sb_sb_0_GPIO_3_M2F                      : out   std_logic;
          DAPI_RX                                 : in    std_logic := 'U';
          DAPI_TX                                 : out   std_logic;
          TM_RX                                   : in    std_logic := 'U';
          TM_TX                                   : out   std_logic
        );
  end component;

  component sb_sb_FABOSC_0_OSC
    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : out   std_logic
        );
  end component;

  component CoreAPB3
    port( sb_sb_0_STAMP_PRDATA                    : in    std_logic_vector(31 downto 0) := (others => 'U');
          sb_sb_0_Memory_PRDATA                   : in    std_logic_vector(31 downto 0) := (others => 'U');
          sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : out   std_logic_vector(31 downto 0);
          STAMP_PADDRS                            : in    std_logic_vector(15 downto 12) := (others => 'U');
          PREADY_N_7                              : out   std_logic;
          sb_sb_0_STAMP_PREADY                    : in    std_logic := 'U';
          sb_sb_0_Memory_PREADY                   : in    std_logic := 'U';
          PRDATA_N_5_i                            : out   std_logic;
          sb_sb_0_STAMP_PSELx                     : out   std_logic;
          sb_sb_0_Memory_PSELx                    : out   std_logic;
          sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx  : in    std_logic := 'U'
        );
  end component;

  component sb_sb_CCC_0_FCCC
    port( FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC : in    std_logic := 'U';
          FIC_0_LOCK                                         : out   std_logic;
          adc_clk_c                                          : out   std_logic;
          sb_sb_0_FIC_0_CLK                                  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \sb_sb_0_FIC_0_CLK\ : std_logic;
    signal sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA : 
        std_logic_vector(31 downto 0);
    signal STAMP_PADDRS : std_logic_vector(15 downto 12);
    signal FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        FIC_0_LOCK, N_2042, PREADY_N_7, PRDATA_N_5_i, 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, N_2043, \GND\, 
        \VCC\ : std_logic;

    for all : sb_sb_MSS
	Use entity work.sb_sb_MSS(DEF_ARCH);
    for all : sb_sb_FABOSC_0_OSC
	Use entity work.sb_sb_FABOSC_0_OSC(DEF_ARCH);
    for all : CoreAPB3
	Use entity work.CoreAPB3(DEF_ARCH);
    for all : sb_sb_CCC_0_FCCC
	Use entity work.sb_sb_CCC_0_FCCC(DEF_ARCH);
begin 

    sb_sb_0_FIC_0_CLK <= \sb_sb_0_FIC_0_CLK\;

    sb_sb_MSS_0 : sb_sb_MSS
      port map(sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(7) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(7), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(6) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(6), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(5) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(5), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(4) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(4), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(3) => N_2043, 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(2) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(2), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(1) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(1), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(0) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(0), dataReady_0
         => dataReady_0, sb_sb_0_STAMP_PWDATA(31) => 
        sb_sb_0_STAMP_PWDATA(31), sb_sb_0_STAMP_PWDATA(30) => 
        sb_sb_0_STAMP_PWDATA(30), sb_sb_0_STAMP_PWDATA(29) => 
        sb_sb_0_STAMP_PWDATA(29), sb_sb_0_STAMP_PWDATA(28) => 
        sb_sb_0_STAMP_PWDATA(28), sb_sb_0_STAMP_PWDATA(27) => 
        sb_sb_0_STAMP_PWDATA(27), sb_sb_0_STAMP_PWDATA(26) => 
        sb_sb_0_STAMP_PWDATA(26), sb_sb_0_STAMP_PWDATA(25) => 
        sb_sb_0_STAMP_PWDATA(25), sb_sb_0_STAMP_PWDATA(24) => 
        sb_sb_0_STAMP_PWDATA(24), sb_sb_0_STAMP_PWDATA(23) => 
        sb_sb_0_STAMP_PWDATA(23), sb_sb_0_STAMP_PWDATA(22) => 
        sb_sb_0_STAMP_PWDATA(22), sb_sb_0_STAMP_PWDATA(21) => 
        sb_sb_0_STAMP_PWDATA(21), sb_sb_0_STAMP_PWDATA(20) => 
        sb_sb_0_STAMP_PWDATA(20), sb_sb_0_STAMP_PWDATA(19) => 
        sb_sb_0_STAMP_PWDATA(19), sb_sb_0_STAMP_PWDATA(18) => 
        sb_sb_0_STAMP_PWDATA(18), sb_sb_0_STAMP_PWDATA(17) => 
        sb_sb_0_STAMP_PWDATA(17), sb_sb_0_STAMP_PWDATA(16) => 
        sb_sb_0_STAMP_PWDATA(16), sb_sb_0_STAMP_PWDATA(15) => 
        sb_sb_0_STAMP_PWDATA(15), sb_sb_0_STAMP_PWDATA(14) => 
        sb_sb_0_STAMP_PWDATA(14), sb_sb_0_STAMP_PWDATA(13) => 
        sb_sb_0_STAMP_PWDATA(13), sb_sb_0_STAMP_PWDATA(12) => 
        sb_sb_0_STAMP_PWDATA(12), sb_sb_0_STAMP_PWDATA(11) => 
        sb_sb_0_STAMP_PWDATA(11), sb_sb_0_STAMP_PWDATA(10) => 
        sb_sb_0_STAMP_PWDATA(10), sb_sb_0_STAMP_PWDATA(9) => 
        sb_sb_0_STAMP_PWDATA(9), sb_sb_0_STAMP_PWDATA(8) => 
        sb_sb_0_STAMP_PWDATA(8), sb_sb_0_STAMP_PWDATA(7) => 
        sb_sb_0_STAMP_PWDATA(7), sb_sb_0_STAMP_PWDATA(6) => 
        sb_sb_0_STAMP_PWDATA(6), sb_sb_0_STAMP_PWDATA(5) => 
        sb_sb_0_STAMP_PWDATA(5), sb_sb_0_STAMP_PWDATA(4) => 
        sb_sb_0_STAMP_PWDATA(4), sb_sb_0_STAMP_PWDATA(3) => 
        sb_sb_0_STAMP_PWDATA(3), sb_sb_0_STAMP_PWDATA(2) => 
        sb_sb_0_STAMP_PWDATA(2), sb_sb_0_STAMP_PWDATA(1) => 
        sb_sb_0_STAMP_PWDATA(1), sb_sb_0_STAMP_PWDATA(0) => 
        sb_sb_0_STAMP_PWDATA(0), STAMP_PADDRS(15) => 
        STAMP_PADDRS(15), STAMP_PADDRS(14) => STAMP_PADDRS(14), 
        STAMP_PADDRS(13) => STAMP_PADDRS(13), STAMP_PADDRS(12)
         => STAMP_PADDRS(12), sb_sb_0_STAMP_PADDR(11) => 
        sb_sb_0_STAMP_PADDR(11), sb_sb_0_STAMP_PADDR(10) => 
        sb_sb_0_STAMP_PADDR(10), sb_sb_0_STAMP_PADDR(9) => 
        sb_sb_0_STAMP_PADDR(9), sb_sb_0_STAMP_PADDR(8) => 
        sb_sb_0_STAMP_PADDR(8), sb_sb_0_STAMP_PADDR(7) => 
        sb_sb_0_STAMP_PADDR(7), sb_sb_0_STAMP_PADDR(6) => 
        sb_sb_0_STAMP_PADDR(6), sb_sb_0_STAMP_PADDR(5) => 
        sb_sb_0_STAMP_PADDR(5), sb_sb_0_STAMP_PADDR(4) => 
        sb_sb_0_STAMP_PADDR(4), sb_sb_0_STAMP_PADDR(3) => 
        sb_sb_0_STAMP_PADDR(3), sb_sb_0_STAMP_PADDR(2) => 
        sb_sb_0_STAMP_PADDR(2), sb_sb_0_STAMP_PADDR(1) => 
        sb_sb_0_STAMP_PADDR(1), sb_sb_0_STAMP_PADDR(0) => 
        sb_sb_0_STAMP_PADDR(0), sb_sb_0_FIC_0_CLK => 
        \sb_sb_0_FIC_0_CLK\, RXSM_SODS_c => RXSM_SODS_c, 
        RXSM_SOE_c => RXSM_SOE_c, RXSM_LO_c => RXSM_LO_c, 
        FIC_0_LOCK => FIC_0_LOCK, PREADY_N_7 => PREADY_N_7, 
        PRDATA_N_5_i => PRDATA_N_5_i, GPIO_6_M2F_c => 
        GPIO_6_M2F_c, LED_RECORDING_c => LED_RECORDING_c, 
        LED_HEARTBEAT_c => LED_HEARTBEAT_c, sb_sb_0_STAMP_PWRITE
         => sb_sb_0_STAMP_PWRITE, 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, 
        sb_sb_0_STAMP_PENABLE => sb_sb_0_STAMP_PENABLE, 
        sb_sb_0_GPIO_4_M2F => sb_sb_0_GPIO_4_M2F, 
        sb_sb_0_GPIO_3_M2F => sb_sb_0_GPIO_3_M2F, DAPI_RX => 
        DAPI_RX, DAPI_TX => DAPI_TX, TM_RX => TM_RX, TM_TX => 
        TM_TX);
    
    FABOSC_0 : sb_sb_FABOSC_0_OSC
      port map(FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
         => FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC);
    
    CoreAPB3_0 : CoreAPB3
      port map(sb_sb_0_STAMP_PRDATA(31) => 
        sb_sb_0_STAMP_PRDATA(31), sb_sb_0_STAMP_PRDATA(30) => 
        sb_sb_0_STAMP_PRDATA(30), sb_sb_0_STAMP_PRDATA(29) => 
        sb_sb_0_STAMP_PRDATA(29), sb_sb_0_STAMP_PRDATA(28) => 
        sb_sb_0_STAMP_PRDATA(28), sb_sb_0_STAMP_PRDATA(27) => 
        sb_sb_0_STAMP_PRDATA(27), sb_sb_0_STAMP_PRDATA(26) => 
        sb_sb_0_STAMP_PRDATA(26), sb_sb_0_STAMP_PRDATA(25) => 
        sb_sb_0_STAMP_PRDATA(25), sb_sb_0_STAMP_PRDATA(24) => 
        sb_sb_0_STAMP_PRDATA(24), sb_sb_0_STAMP_PRDATA(23) => 
        sb_sb_0_STAMP_PRDATA(23), sb_sb_0_STAMP_PRDATA(22) => 
        sb_sb_0_STAMP_PRDATA(22), sb_sb_0_STAMP_PRDATA(21) => 
        sb_sb_0_STAMP_PRDATA(21), sb_sb_0_STAMP_PRDATA(20) => 
        sb_sb_0_STAMP_PRDATA(20), sb_sb_0_STAMP_PRDATA(19) => 
        sb_sb_0_STAMP_PRDATA(19), sb_sb_0_STAMP_PRDATA(18) => 
        sb_sb_0_STAMP_PRDATA(18), sb_sb_0_STAMP_PRDATA(17) => 
        sb_sb_0_STAMP_PRDATA(17), sb_sb_0_STAMP_PRDATA(16) => 
        sb_sb_0_STAMP_PRDATA(16), sb_sb_0_STAMP_PRDATA(15) => 
        sb_sb_0_STAMP_PRDATA(15), sb_sb_0_STAMP_PRDATA(14) => 
        sb_sb_0_STAMP_PRDATA(14), sb_sb_0_STAMP_PRDATA(13) => 
        sb_sb_0_STAMP_PRDATA(13), sb_sb_0_STAMP_PRDATA(12) => 
        sb_sb_0_STAMP_PRDATA(12), sb_sb_0_STAMP_PRDATA(11) => 
        sb_sb_0_STAMP_PRDATA(11), sb_sb_0_STAMP_PRDATA(10) => 
        sb_sb_0_STAMP_PRDATA(10), sb_sb_0_STAMP_PRDATA(9) => 
        sb_sb_0_STAMP_PRDATA(9), sb_sb_0_STAMP_PRDATA(8) => 
        sb_sb_0_STAMP_PRDATA(8), sb_sb_0_STAMP_PRDATA(7) => 
        sb_sb_0_STAMP_PRDATA(7), sb_sb_0_STAMP_PRDATA(6) => 
        sb_sb_0_STAMP_PRDATA(6), sb_sb_0_STAMP_PRDATA(5) => 
        sb_sb_0_STAMP_PRDATA(5), sb_sb_0_STAMP_PRDATA(4) => 
        sb_sb_0_STAMP_PRDATA(4), sb_sb_0_STAMP_PRDATA(3) => 
        sb_sb_0_STAMP_PRDATA(3), sb_sb_0_STAMP_PRDATA(2) => 
        sb_sb_0_STAMP_PRDATA(2), sb_sb_0_STAMP_PRDATA(1) => 
        sb_sb_0_STAMP_PRDATA(1), sb_sb_0_STAMP_PRDATA(0) => 
        sb_sb_0_STAMP_PRDATA(0), sb_sb_0_Memory_PRDATA(31) => 
        sb_sb_0_Memory_PRDATA(31), sb_sb_0_Memory_PRDATA(30) => 
        sb_sb_0_Memory_PRDATA(30), sb_sb_0_Memory_PRDATA(29) => 
        sb_sb_0_Memory_PRDATA(29), sb_sb_0_Memory_PRDATA(28) => 
        sb_sb_0_Memory_PRDATA(28), sb_sb_0_Memory_PRDATA(27) => 
        sb_sb_0_Memory_PRDATA(27), sb_sb_0_Memory_PRDATA(26) => 
        sb_sb_0_Memory_PRDATA(26), sb_sb_0_Memory_PRDATA(25) => 
        sb_sb_0_Memory_PRDATA(25), sb_sb_0_Memory_PRDATA(24) => 
        sb_sb_0_Memory_PRDATA(24), sb_sb_0_Memory_PRDATA(23) => 
        sb_sb_0_Memory_PRDATA(23), sb_sb_0_Memory_PRDATA(22) => 
        sb_sb_0_Memory_PRDATA(22), sb_sb_0_Memory_PRDATA(21) => 
        sb_sb_0_Memory_PRDATA(21), sb_sb_0_Memory_PRDATA(20) => 
        sb_sb_0_Memory_PRDATA(20), sb_sb_0_Memory_PRDATA(19) => 
        sb_sb_0_Memory_PRDATA(19), sb_sb_0_Memory_PRDATA(18) => 
        sb_sb_0_Memory_PRDATA(18), sb_sb_0_Memory_PRDATA(17) => 
        sb_sb_0_Memory_PRDATA(17), sb_sb_0_Memory_PRDATA(16) => 
        sb_sb_0_Memory_PRDATA(16), sb_sb_0_Memory_PRDATA(15) => 
        sb_sb_0_Memory_PRDATA(15), sb_sb_0_Memory_PRDATA(14) => 
        sb_sb_0_Memory_PRDATA(14), sb_sb_0_Memory_PRDATA(13) => 
        sb_sb_0_Memory_PRDATA(13), sb_sb_0_Memory_PRDATA(12) => 
        sb_sb_0_Memory_PRDATA(12), sb_sb_0_Memory_PRDATA(11) => 
        sb_sb_0_Memory_PRDATA(11), sb_sb_0_Memory_PRDATA(10) => 
        sb_sb_0_Memory_PRDATA(10), sb_sb_0_Memory_PRDATA(9) => 
        sb_sb_0_Memory_PRDATA(9), sb_sb_0_Memory_PRDATA(8) => 
        sb_sb_0_Memory_PRDATA(8), sb_sb_0_Memory_PRDATA(7) => 
        sb_sb_0_Memory_PRDATA(7), sb_sb_0_Memory_PRDATA(6) => 
        sb_sb_0_Memory_PRDATA(6), sb_sb_0_Memory_PRDATA(5) => 
        sb_sb_0_Memory_PRDATA(5), sb_sb_0_Memory_PRDATA(4) => 
        sb_sb_0_Memory_PRDATA(4), sb_sb_0_Memory_PRDATA(3) => 
        sb_sb_0_Memory_PRDATA(3), sb_sb_0_Memory_PRDATA(2) => 
        sb_sb_0_Memory_PRDATA(2), sb_sb_0_Memory_PRDATA(1) => 
        sb_sb_0_Memory_PRDATA(1), sb_sb_0_Memory_PRDATA(0) => 
        sb_sb_0_Memory_PRDATA(0), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(31), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(30), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(29), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(28), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(27), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(26), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(25), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(24), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(23), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(22), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(21), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(20), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(19), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(18), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(17), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(16), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(15), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(14), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(13), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(12), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(11), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(10), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(9), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(8), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(7) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(7), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(6) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(6), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(5) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(5), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(4) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(4), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(3) => N_2042, 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(2) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(2), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(1) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(1), 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(0) => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA(0), 
        STAMP_PADDRS(15) => STAMP_PADDRS(15), STAMP_PADDRS(14)
         => STAMP_PADDRS(14), STAMP_PADDRS(13) => 
        STAMP_PADDRS(13), STAMP_PADDRS(12) => STAMP_PADDRS(12), 
        PREADY_N_7 => PREADY_N_7, sb_sb_0_STAMP_PREADY => 
        sb_sb_0_STAMP_PREADY, sb_sb_0_Memory_PREADY => 
        sb_sb_0_Memory_PREADY, PRDATA_N_5_i => PRDATA_N_5_i, 
        sb_sb_0_STAMP_PSELx => sb_sb_0_STAMP_PSELx, 
        sb_sb_0_Memory_PSELx => sb_sb_0_Memory_PSELx, 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx => 
        sb_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx);
    
    CCC_0 : sb_sb_CCC_0_FCCC
      port map(FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
         => FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        FIC_0_LOCK => FIC_0_LOCK, adc_clk_c => adc_clk_c, 
        sb_sb_0_FIC_0_CLK => \sb_sb_0_FIC_0_CLK\);
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => sb_sb_0_POWER_ON_RESET_N, 
        DEVRST_N => DEVRST_N);
    
    GND_Z : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity spi_master_1_16 is

    port( component_state_0      : in    std_logic;
          spi_tx_data            : in    std_logic_vector(15 downto 0);
          spi_rx_data            : out   std_logic_vector(15 downto 0);
          delay_countere         : out   std_logic;
          N_176                  : in    std_logic;
          delay_counterlde_0_0_0 : in    std_logic;
          enable                 : in    std_logic;
          spi_busy               : out   std_logic;
          mosi_cl_0              : out   std_logic;
          mosi_1_0               : out   std_logic;
          debug_led_net_0        : in    std_logic;
          stamp0_spi_clock_c     : out   std_logic;
          debug_led_net_0_arst   : in    std_logic;
          stamp0_spi_miso_c      : in    std_logic;
          sb_sb_0_FIC_0_CLK      : in    std_logic
        );

end spi_master_1_16;

architecture DEF_ARCH of spi_master_1_16 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \spi_busy\, \mosi_cl_0\, \stamp0_spi_clock_c\
         : std_logic;
    signal rx_buffer_Z : std_logic_vector(15 downto 0);
    signal tx_buffer_Z : std_logic_vector(15 downto 0);
    signal ss_n_buffer_Z : std_logic_vector(0 to 0);
    signal state_Z : std_logic_vector(0 to 0);
    signal clk_toggles_Z : std_logic_vector(5 downto 0);
    signal clk_toggles_lm : std_logic_vector(5 downto 0);
    signal count_Z : std_logic_vector(31 downto 0);
    signal count_lm : std_logic_vector(31 downto 0);
    signal count_cry_Z : std_logic_vector(30 downto 1);
    signal count_s : std_logic_vector(30 downto 1);
    signal count_cry_Y : std_logic_vector(30 downto 1);
    signal count_s_FCO : std_logic_vector(31 to 31);
    signal count_s_Z : std_logic_vector(31 to 31);
    signal count_s_Y : std_logic_vector(31 to 31);
    signal clk_toggles_cry_Z : std_logic_vector(4 downto 1);
    signal clk_toggles_s : std_logic_vector(4 downto 1);
    signal clk_toggles_cry_Y : std_logic_vector(4 downto 1);
    signal clk_toggles_s_FCO : std_logic_vector(5 to 5);
    signal clk_toggles_s_Z : std_logic_vector(5 to 5);
    signal clk_toggles_s_Y : std_logic_vector(5 to 5);
    signal \VCC\, rx_buffer_0_sqmuxa_1, \GND\, N_219, 
        un1_reset_n_inv_2_i, N_218, N_217, N_216, N_215, N_214, 
        N_213, N_212, N_211, N_210, N_209, N_208, N_207, N_206, 
        N_205, N_50_i, N_333, N_20_i, assert_data_Z, N_186_i, 
        mosi_1_1, N_192, busy_7, N_25_i, N_37_i, N_49_i, 
        count_s_832_FCO, count_s_832_S, count_s_832_Y, 
        clk_toggles_s_833_FCO, clk_toggles_s_833_S, 
        clk_toggles_s_833_Y, un7_count_NE_i, 
        un1_reset_n_inv_2_i_1, N_322, 
        rx_buffer_0_sqmuxa_1_0_a2_3_a3_0_Z, un7_count_NE_13_Z, 
        N_320, un7_count_NE_23_Z, un7_count_NE_21_Z, 
        un7_count_NE_20_Z, un7_count_NE_19_Z, un7_count_NE_18_Z, 
        un7_count_NE_17_Z, un7_count_NE_16_Z, 
        un10_count_0_a2_0_a3_3_Z, 
        rx_buffer_0_sqmuxa_1_0_a2_3_a2_2_Z, count_0_sqmuxa, 
        un10_count_i, un7_count_NE_27_Z, mosi_cl_4_i_0_1_Z, 
        un7_count_NE_28_Z, N_312, sclk_buffer_0_sqmuxa, N_1489, 
        N_68 : std_logic;

begin 

    spi_busy <= \spi_busy\;
    mosi_cl_0 <= \mosi_cl_0\;
    stamp0_spi_clock_c <= \stamp0_spi_clock_c\;

    \count_lm_0[13]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(13), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(13));
    
    \count[27]\ : SLE
      port map(D => count_lm(27), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(27));
    
    \rx_buffer[11]\ : SLE
      port map(D => rx_buffer_Z(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(11));
    
    \state[0]\ : SLE
      port map(D => busy_7, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => state_Z(0));
    
    \count[25]\ : SLE
      port map(D => count_lm(25), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(25));
    
    \tx_buffer_RNO[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(14), B => tx_buffer_Z(13), C => 
        state_Z(0), Y => N_206);
    
    \count[17]\ : SLE
      port map(D => count_lm(17), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(17));
    
    \tx_buffer[11]\ : SLE
      port map(D => N_209, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(11));
    
    \count[15]\ : SLE
      port map(D => count_lm(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(15));
    
    \count_cry[14]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(14), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(13), S => count_s(14), Y => 
        count_cry_Y(14), FCO => count_cry_Z(14));
    
    \rx_data[2]\ : SLE
      port map(D => rx_buffer_Z(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(2));
    
    \count[9]\ : SLE
      port map(D => count_lm(9), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(9));
    
    \state_RNIDMJE[0]\ : CFG3
      generic map(INIT => x"E0")

      port map(A => enable, B => state_Z(0), C => debug_led_net_0, 
        Y => N_49_i);
    
    \count_lm_0[17]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(17), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(17));
    
    \count_cry[28]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(28), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(27), S => count_s(28), Y => 
        count_cry_Y(28), FCO => count_cry_Z(28));
    
    \count[8]\ : SLE
      port map(D => count_lm(8), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(8));
    
    \count_cry[26]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(26), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(25), S => count_s(26), Y => 
        count_cry_Y(26), FCO => count_cry_Z(26));
    
    \clk_toggles_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => clk_toggles_Z(2), C => \GND\, D
         => \GND\, FCI => clk_toggles_cry_Z(1), S => 
        clk_toggles_s(2), Y => clk_toggles_cry_Y(2), FCO => 
        clk_toggles_cry_Z(2));
    
    \rx_data[15]\ : SLE
      port map(D => rx_buffer_Z(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(15));
    
    \count_cry[20]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(20), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(19), S => count_s(20), Y => 
        count_cry_Y(20), FCO => count_cry_Z(20));
    
    \count_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(8), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(7), S => count_s(8), Y => 
        count_cry_Y(8), FCO => count_cry_Z(8));
    
    \count_lm_0[6]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(6), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(6));
    
    \rx_data[3]\ : SLE
      port map(D => rx_buffer_Z(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(3));
    
    \rx_data[7]\ : SLE
      port map(D => rx_buffer_Z(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(7));
    
    \tx_buffer[5]\ : SLE
      port map(D => N_215, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(5));
    
    \tx_buffer_RNO[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(1), B => tx_buffer_Z(0), C => 
        state_Z(0), Y => N_219);
    
    \tx_buffer_RNO[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(13), B => tx_buffer_Z(12), C => 
        state_Z(0), Y => N_207);
    
    rx_buffer_0_sqmuxa_1_0_a2_3_a2_2 : CFG3
      generic map(INIT => x"01")

      port map(A => clk_toggles_Z(3), B => clk_toggles_Z(1), C
         => clk_toggles_Z(0), Y => 
        rx_buffer_0_sqmuxa_1_0_a2_3_a2_2_Z);
    
    \rx_buffer[10]\ : SLE
      port map(D => rx_buffer_Z(9), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(10));
    
    \count[20]\ : SLE
      port map(D => count_lm(20), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(20));
    
    \rx_data[4]\ : SLE
      port map(D => rx_buffer_Z(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(4));
    
    \tx_buffer[10]\ : SLE
      port map(D => N_210, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(10));
    
    \count_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(2), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(1), S => count_s(2), Y => 
        count_cry_Y(2), FCO => count_cry_Z(2));
    
    \count[10]\ : SLE
      port map(D => count_lm(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(10));
    
    \tx_buffer[7]\ : SLE
      port map(D => N_213, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(7));
    
    \tx_buffer[3]\ : SLE
      port map(D => N_217, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(3));
    
    \count_lm_0[5]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(5), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(5));
    
    \count_lm_0[28]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(28), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(28));
    
    \count_cry[15]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(15), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(14), S => count_s(15), Y => 
        count_cry_Y(15), FCO => count_cry_Z(15));
    
    \clk_toggles_lm_0[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_192, B => clk_toggles_Z(0), Y => 
        clk_toggles_lm(0));
    
    \count[5]\ : SLE
      port map(D => count_lm(5), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(5));
    
    \rx_buffer[14]\ : SLE
      port map(D => rx_buffer_Z(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(14));
    
    \clk_toggles_lm_0[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_192, B => clk_toggles_s_Z(5), Y => 
        clk_toggles_lm(5));
    
    un10_count_0_a2_0_a3 : CFG3
      generic map(INIT => x"80")

      port map(A => clk_toggles_Z(0), B => 
        un10_count_0_a2_0_a3_3_Z, C => clk_toggles_Z(5), Y => 
        un10_count_i);
    
    \tx_buffer_RNO[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(9), B => tx_buffer_Z(8), C => 
        state_Z(0), Y => N_211);
    
    \count_s[31]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(31), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(30), S => count_s_Z(31), Y => 
        count_s_Y(31), FCO => count_s_FCO(31));
    
    \tx_buffer_RNO[6]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(6), B => tx_buffer_Z(5), C => 
        state_Z(0), Y => N_214);
    
    \tx_buffer[14]\ : SLE
      port map(D => N_206, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(14));
    
    \rx_data[5]\ : SLE
      port map(D => rx_buffer_Z(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(5));
    
    \rx_buffer[7]\ : SLE
      port map(D => rx_buffer_Z(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(7));
    
    \rx_buffer[13]\ : SLE
      port map(D => rx_buffer_Z(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(13));
    
    un7_count_NE_16 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(7), B => count_Z(6), C => count_Z(5), 
        D => count_Z(4), Y => un7_count_NE_16_Z);
    
    \tx_buffer_RNO[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(15), B => tx_buffer_Z(14), C => 
        state_Z(0), Y => N_205);
    
    \count_cry[30]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(30), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(29), S => count_s(30), Y => 
        count_cry_Y(30), FCO => count_cry_Z(30));
    
    \count_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(12), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(11), S => count_s(12), Y => 
        count_cry_Y(12), FCO => count_cry_Z(12));
    
    \tx_buffer[13]\ : SLE
      port map(D => N_207, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(13));
    
    \count_lm_0[24]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(24), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(24));
    
    \count_cry[19]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(19), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(18), S => count_s(19), Y => 
        count_cry_Y(19), FCO => count_cry_Z(19));
    
    \count[4]\ : SLE
      port map(D => count_lm(4), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(4));
    
    \clk_toggles_lm_0[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_192, B => clk_toggles_s(2), Y => 
        clk_toggles_lm(2));
    
    sclk_buffer_RNO : CFG4
      generic map(INIT => x"2788")

      port map(A => state_Z(0), B => sclk_buffer_0_sqmuxa, C => 
        enable, D => \stamp0_spi_clock_c\, Y => N_20_i);
    
    \count[22]\ : SLE
      port map(D => count_lm(22), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(22));
    
    mosi_1 : SLE
      port map(D => tx_buffer_Z(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => mosi_1_1, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => mosi_1_0);
    
    \count[12]\ : SLE
      port map(D => count_lm(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(12));
    
    \count_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(6), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(5), S => count_s(6), Y => 
        count_cry_Y(6), FCO => count_cry_Z(6));
    
    \count[0]\ : SLE
      port map(D => count_lm(0), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(0));
    
    assert_data_RNO : CFG4
      generic map(INIT => x"82C3")

      port map(A => state_Z(0), B => N_320, C => assert_data_Z, D
         => enable, Y => N_186_i);
    
    \rx_data[11]\ : SLE
      port map(D => rx_buffer_Z(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(11));
    
    \count_lm_0[21]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(21), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(21));
    
    mosi_cl_4_i_0_o2_RNIIPO72 : CFG4
      generic map(INIT => x"4030")

      port map(A => N_322, B => state_Z(0), C => debug_led_net_0, 
        D => un1_reset_n_inv_2_i_1, Y => un1_reset_n_inv_2_i);
    
    \count_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(5), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(4), S => count_s(5), Y => 
        count_cry_Y(5), FCO => count_cry_Z(5));
    
    \tx_buffer_RNO[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(2), B => tx_buffer_Z(1), C => 
        state_Z(0), Y => N_218);
    
    \rx_buffer[8]\ : SLE
      port map(D => rx_buffer_Z(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(8));
    
    rx_buffer_0_sqmuxa_1_0_a2_3_o2 : CFG4
      generic map(INIT => x"10FF")

      port map(A => clk_toggles_Z(2), B => clk_toggles_Z(4), C
         => rx_buffer_0_sqmuxa_1_0_a2_3_a2_2_Z, D => 
        clk_toggles_Z(5), Y => N_312);
    
    \tx_buffer[9]\ : SLE
      port map(D => N_211, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(9));
    
    \count_lm_0[8]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(8), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(8));
    
    \tx_buffer_RNO[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(4), B => tx_buffer_Z(3), C => 
        state_Z(0), Y => N_216);
    
    \tx_buffer[2]\ : SLE
      port map(D => N_218, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(2));
    
    \count_lm_0[10]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(10), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(10));
    
    \rx_buffer[5]\ : SLE
      port map(D => rx_buffer_Z(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(5));
    
    \count_lm_0[29]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(29), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(29));
    
    \clk_toggles_lm_0[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_192, B => clk_toggles_s(4), Y => 
        clk_toggles_lm(4));
    
    \rx_buffer[4]\ : SLE
      port map(D => rx_buffer_Z(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(4));
    
    \count_cry[21]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(21), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(20), S => count_s(21), Y => 
        count_cry_Y(21), FCO => count_cry_Z(21));
    
    count_s_832 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(0), C => \GND\, D => 
        \GND\, FCI => \VCC\, S => count_s_832_S, Y => 
        count_s_832_Y, FCO => count_s_832_FCO);
    
    \count[23]\ : SLE
      port map(D => count_lm(23), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(23));
    
    busy : SLE
      port map(D => busy_7, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => debug_led_net_0_arst, ADn => \GND\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => \spi_busy\);
    
    \count[13]\ : SLE
      port map(D => count_lm(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(13));
    
    \count_cry[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(13), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(12), S => count_s(13), Y => 
        count_cry_Y(13), FCO => count_cry_Z(13));
    
    \count_cry[24]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(24), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(23), S => count_s(24), Y => 
        count_cry_Y(24), FCO => count_cry_Z(24));
    
    mosi_cl_4_i_0_o2 : CFG2
      generic map(INIT => x"B")

      port map(A => clk_toggles_Z(5), B => assert_data_Z, Y => 
        N_322);
    
    \state_RNID0SF1[0]\ : CFG3
      generic map(INIT => x"8D")

      port map(A => state_Z(0), B => un7_count_NE_i, C => enable, 
        Y => un1_reset_n_inv_2_i_1);
    
    \count_cry[17]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(17), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(16), S => count_s(17), Y => 
        count_cry_Y(17), FCO => count_cry_Z(17));
    
    GND_Z : GND
      port map(Y => \GND\);
    
    un7_count_NE_17 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(11), B => count_Z(10), C => 
        count_Z(9), D => count_Z(8), Y => un7_count_NE_17_Z);
    
    un7_count_NE_18 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(15), B => count_Z(14), C => 
        count_Z(13), D => count_Z(12), Y => un7_count_NE_18_Z);
    
    \clk_toggles_lm_0[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_192, B => clk_toggles_s(3), Y => 
        clk_toggles_lm(3));
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    un10_count_0_a2_0_a3_RNIF61H : CFG2
      generic map(INIT => x"4")

      port map(A => N_320, B => un10_count_i, Y => N_50_i);
    
    ss_n_buffer_1_sqmuxa_0_a2_i : CFG3
      generic map(INIT => x"B3")

      port map(A => un7_count_NE_i, B => state_Z(0), C => 
        un10_count_i, Y => N_192);
    
    \count_lm_0[0]\ : CFG3
      generic map(INIT => x"F7")

      port map(A => count_Z(0), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(0));
    
    \count_lm_0[25]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(25), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(25));
    
    un7_count_NE_13 : CFG2
      generic map(INIT => x"E")

      port map(A => count_Z(30), B => count_Z(31), Y => 
        un7_count_NE_13_Z);
    
    \rx_data[1]\ : SLE
      port map(D => rx_buffer_Z(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(1));
    
    \rx_buffer[1]\ : SLE
      port map(D => rx_buffer_Z(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(1));
    
    \rx_data[14]\ : SLE
      port map(D => rx_buffer_Z(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(14));
    
    \count[1]\ : SLE
      port map(D => count_lm(1), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(1));
    
    \count[3]\ : SLE
      port map(D => count_lm(3), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(3));
    
    busy_RNI9S1EA : CFG4
      generic map(INIT => x"F0FD")

      port map(A => \spi_busy\, B => component_state_0, C => 
        delay_counterlde_0_0_0, D => N_176, Y => delay_countere);
    
    \rx_buffer[15]\ : SLE
      port map(D => rx_buffer_Z(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(15));
    
    \clk_toggles[2]\ : SLE
      port map(D => clk_toggles_lm(2), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_37_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => clk_toggles_Z(2));
    
    \rx_buffer[12]\ : SLE
      port map(D => rx_buffer_Z(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(12));
    
    \count_lm_0[4]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(4), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(4));
    
    \count_lm_0[22]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(22), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(22));
    
    \count[29]\ : SLE
      port map(D => count_lm(29), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(29));
    
    \count_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(7), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(6), S => count_s(7), Y => 
        count_cry_Y(7), FCO => count_cry_Z(7));
    
    \tx_buffer[15]\ : SLE
      port map(D => N_205, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(15));
    
    \count[19]\ : SLE
      port map(D => count_lm(19), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(19));
    
    \tx_buffer[12]\ : SLE
      port map(D => N_208, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(12));
    
    \count_lm_0[18]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(18), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(18));
    
    un7_count_NE_27 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(28), B => count_Z(29), C => 
        un7_count_NE_23_Z, D => un7_count_NE_13_Z, Y => 
        un7_count_NE_27_Z);
    
    un7_count_NE_28 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un7_count_NE_19_Z, B => un7_count_NE_18_Z, C
         => un7_count_NE_17_Z, D => un7_count_NE_16_Z, Y => 
        un7_count_NE_28_Z);
    
    \clk_toggles[0]\ : SLE
      port map(D => clk_toggles_lm(0), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_37_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => clk_toggles_Z(0));
    
    \tx_buffer[4]\ : SLE
      port map(D => N_216, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(4));
    
    \count_lm_0[30]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(30), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(30));
    
    un7_count_NE_23 : CFG4
      generic map(INIT => x"7FFF")

      port map(A => count_Z(3), B => count_Z(2), C => count_Z(1), 
        D => count_Z(0), Y => un7_count_NE_23_Z);
    
    \count_cry[25]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(25), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(24), S => count_s(25), Y => 
        count_cry_Y(25), FCO => count_cry_Z(25));
    
    \clk_toggles[1]\ : SLE
      port map(D => clk_toggles_lm(1), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_37_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => clk_toggles_Z(1));
    
    mosi_cl_4_i_0_1 : CFG4
      generic map(INIT => x"7F5F")

      port map(A => state_Z(0), B => \mosi_cl_0\, C => 
        debug_led_net_0, D => N_322, Y => mosi_cl_4_i_0_1_Z);
    
    sclk_buffer : SLE
      port map(D => N_20_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        debug_led_net_0, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => \stamp0_spi_clock_c\);
    
    \count_lm_0[26]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(26), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(26));
    
    \count_lm_0[9]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(9), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(9));
    
    \rx_buffer[3]\ : SLE
      port map(D => rx_buffer_Z(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(3));
    
    \tx_buffer[8]\ : SLE
      port map(D => N_212, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(8));
    
    \count_lm_0[14]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(14), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(14));
    
    un7_count_NE_19 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(19), B => count_Z(18), C => 
        count_Z(17), D => count_Z(16), Y => un7_count_NE_19_Z);
    
    rx_data_0_sqmuxa_i_0_o3_RNIHNAO : CFG4
      generic map(INIT => x"44C4")

      port map(A => N_320, B => debug_led_net_0, C => enable, D
         => state_Z(0), Y => N_37_i);
    
    \tx_buffer[6]\ : SLE
      port map(D => N_214, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(6));
    
    \count_cry[22]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(22), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(21), S => count_s(22), Y => 
        count_cry_Y(22), FCO => count_cry_Z(22));
    
    \count_cry[29]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(29), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(28), S => count_s(29), Y => 
        count_cry_Y(29), FCO => count_cry_Z(29));
    
    \tx_buffer_RNO[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => state_Z(0), B => spi_tx_data(0), Y => N_333);
    
    busy_7_0_0_0 : CFG4
      generic map(INIT => x"DDC0")

      port map(A => un10_count_i, B => N_320, C => enable, D => 
        state_Z(0), Y => busy_7);
    
    un7_count_NE_20 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(23), B => count_Z(22), C => 
        count_Z(21), D => count_Z(20), Y => un7_count_NE_20_Z);
    
    \tx_buffer_RNO[5]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(5), B => tx_buffer_Z(4), C => 
        state_Z(0), Y => N_215);
    
    \count_lm_0[23]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(23), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(23));
    
    \count_lm_0[1]\ : CFG4
      generic map(INIT => x"D8CC")

      port map(A => un7_count_NE_i, B => count_0_sqmuxa, C => 
        count_s(1), D => state_Z(0), Y => count_lm(1));
    
    \rx_buffer[6]\ : SLE
      port map(D => rx_buffer_Z(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(6));
    
    \clk_toggles[4]\ : SLE
      port map(D => clk_toggles_lm(4), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_37_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => clk_toggles_Z(4));
    
    mosi_1_1_0_a2_0_a3 : CFG4
      generic map(INIT => x"0004")

      port map(A => N_320, B => debug_led_net_0, C => N_322, D
         => un10_count_i, Y => mosi_1_1);
    
    \count_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(4), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(3), S => count_s(4), Y => 
        count_cry_Y(4), FCO => count_cry_Z(4));
    
    count_0_sqmuxa_0_a2_0_a3 : CFG3
      generic map(INIT => x"20")

      port map(A => enable, B => state_Z(0), C => debug_led_net_0, 
        Y => count_0_sqmuxa);
    
    \count_lm_0[11]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(11), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(11));
    
    \count_cry[18]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(18), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(17), S => count_s(18), Y => 
        count_cry_Y(18), FCO => count_cry_Z(18));
    
    \count_lm_0[27]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s(27), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(27));
    
    \count_cry[16]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(16), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(15), S => count_s(16), Y => 
        count_cry_Y(16), FCO => count_cry_Z(16));
    
    \tx_buffer[1]\ : SLE
      port map(D => N_219, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(1));
    
    \rx_buffer[2]\ : SLE
      port map(D => rx_buffer_Z(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(2));
    
    \count_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(10), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(9), S => count_s(10), Y => 
        count_cry_Y(10), FCO => count_cry_Z(10));
    
    \tx_buffer_RNO[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(12), B => tx_buffer_Z(11), C => 
        state_Z(0), Y => N_208);
    
    \rx_data[10]\ : SLE
      port map(D => rx_buffer_Z(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(10));
    
    \rx_data[12]\ : SLE
      port map(D => rx_buffer_Z(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(12));
    
    \count[31]\ : SLE
      port map(D => count_lm(31), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(31));
    
    \count[28]\ : SLE
      port map(D => count_lm(28), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(28));
    
    \count_lm_0[19]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(19), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(19));
    
    \count[18]\ : SLE
      port map(D => count_lm(18), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(18));
    
    \count[7]\ : SLE
      port map(D => count_lm(7), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(7));
    
    \count_lm_0[3]\ : CFG4
      generic map(INIT => x"D8CC")

      port map(A => un7_count_NE_i, B => count_0_sqmuxa, C => 
        count_s(3), D => state_Z(0), Y => count_lm(3));
    
    \tx_buffer_RNO[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(10), B => tx_buffer_Z(9), C => 
        state_Z(0), Y => N_210);
    
    \clk_toggles_lm_0[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_192, B => clk_toggles_s(1), Y => 
        clk_toggles_lm(1));
    
    un10_count_0_a2_0_a3_3 : CFG4
      generic map(INIT => x"0001")

      port map(A => clk_toggles_Z(4), B => clk_toggles_Z(3), C
         => clk_toggles_Z(2), D => clk_toggles_Z(1), Y => 
        un10_count_0_a2_0_a3_3_Z);
    
    \clk_toggles_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => clk_toggles_Z(1), C => \GND\, D
         => \GND\, FCI => clk_toggles_s_833_FCO, S => 
        clk_toggles_s(1), Y => clk_toggles_cry_Y(1), FCO => 
        clk_toggles_cry_Z(1));
    
    \rx_buffer[0]\ : SLE
      port map(D => stamp0_spi_miso_c, CLK => sb_sb_0_FIC_0_CLK, 
        EN => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        rx_buffer_Z(0));
    
    \rx_buffer[9]\ : SLE
      port map(D => rx_buffer_Z(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => rx_buffer_0_sqmuxa_1, ALn => \VCC\, ADn => \VCC\, SLn
         => \VCC\, SD => \GND\, LAT => \GND\, Q => rx_buffer_Z(9));
    
    \rx_data[8]\ : SLE
      port map(D => rx_buffer_Z(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(8));
    
    \count[6]\ : SLE
      port map(D => count_lm(6), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(6));
    
    \rx_data[6]\ : SLE
      port map(D => rx_buffer_Z(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(6));
    
    clk_toggles_s_833 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => clk_toggles_Z(0), C => \GND\, D
         => \GND\, FCI => \VCC\, S => clk_toggles_s_833_S, Y => 
        clk_toggles_s_833_Y, FCO => clk_toggles_s_833_FCO);
    
    \count_cry[23]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(23), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(22), S => count_s(23), Y => 
        count_cry_Y(23), FCO => count_cry_Z(23));
    
    rx_buffer_0_sqmuxa_1_0_a2_3_a3_0 : CFG2
      generic map(INIT => x"1")

      port map(A => assert_data_Z, B => ss_n_buffer_Z(0), Y => 
        rx_buffer_0_sqmuxa_1_0_a2_3_a3_0_Z);
    
    \ss_n_buffer[0]\ : SLE
      port map(D => N_192, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => debug_led_net_0_arst, ADn => \GND\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => ss_n_buffer_Z(0));
    
    \count_cry[27]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(27), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(26), S => count_s(27), Y => 
        count_cry_Y(27), FCO => count_cry_Z(27));
    
    \count_lm_0[15]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(15), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(15));
    
    \clk_toggles_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => clk_toggles_Z(4), C => \GND\, D
         => \GND\, FCI => clk_toggles_cry_Z(3), S => 
        clk_toggles_s(4), Y => clk_toggles_cry_Y(4), FCO => 
        clk_toggles_cry_Z(4));
    
    \rx_data[0]\ : SLE
      port map(D => rx_buffer_Z(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(0));
    
    rx_buffer_0_sqmuxa_1_0_a2_3_a3 : CFG4
      generic map(INIT => x"0080")

      port map(A => N_312, B => 
        rx_buffer_0_sqmuxa_1_0_a2_3_a3_0_Z, C => debug_led_net_0, 
        D => N_320, Y => rx_buffer_0_sqmuxa_1);
    
    \count[26]\ : SLE
      port map(D => count_lm(26), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(26));
    
    \tx_buffer[0]\ : SLE
      port map(D => N_333, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_reset_n_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => tx_buffer_Z(0));
    
    \count[16]\ : SLE
      port map(D => count_lm(16), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(16));
    
    sclk_buffer_0_sqmuxa_0_a2_0_a3 : CFG3
      generic map(INIT => x"08")

      port map(A => N_312, B => un7_count_NE_i, C => 
        ss_n_buffer_Z(0), Y => sclk_buffer_0_sqmuxa);
    
    \count_lm_0[31]\ : CFG3
      generic map(INIT => x"20")

      port map(A => count_s_Z(31), B => un7_count_NE_i, C => 
        state_Z(0), Y => count_lm(31));
    
    \tx_buffer_RNO[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(8), B => tx_buffer_Z(7), C => 
        state_Z(0), Y => N_212);
    
    \count_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(3), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(2), S => count_s(3), Y => 
        count_cry_Y(3), FCO => count_cry_Z(3));
    
    \count[2]\ : SLE
      port map(D => count_lm(2), CLK => sb_sb_0_FIC_0_CLK, EN => 
        N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => count_Z(2));
    
    \clk_toggles[5]\ : SLE
      port map(D => clk_toggles_lm(5), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_37_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => clk_toggles_Z(5));
    
    \count_lm_0[12]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(12), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(12));
    
    un7_count_NE_20_RNIK2531 : CFG4
      generic map(INIT => x"0001")

      port map(A => un7_count_NE_21_Z, B => un7_count_NE_20_Z, C
         => un7_count_NE_28_Z, D => un7_count_NE_27_Z, Y => 
        un7_count_NE_i);
    
    \clk_toggles[3]\ : SLE
      port map(D => clk_toggles_lm(3), CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_37_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => clk_toggles_Z(3));
    
    un7_count_NE_21 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => count_Z(27), B => count_Z(26), C => 
        count_Z(25), D => count_Z(24), Y => un7_count_NE_21_Z);
    
    \rx_data[13]\ : SLE
      port map(D => rx_buffer_Z(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(13));
    
    \clk_toggles_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => clk_toggles_Z(3), C => \GND\, D
         => \GND\, FCI => clk_toggles_cry_Z(2), S => 
        clk_toggles_s(3), Y => clk_toggles_cry_Y(3), FCO => 
        clk_toggles_cry_Z(3));
    
    \count[21]\ : SLE
      port map(D => count_lm(21), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(21));
    
    mosi_cl : SLE
      port map(D => N_25_i, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => \mosi_cl_0\);
    
    \count[11]\ : SLE
      port map(D => count_lm(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(11));
    
    \clk_toggles_s[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => clk_toggles_Z(5), C => \GND\, D
         => \GND\, FCI => clk_toggles_cry_Z(4), S => 
        clk_toggles_s_Z(5), Y => clk_toggles_s_Y(5), FCO => 
        clk_toggles_s_FCO(5));
    
    \count_lm_0[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(7), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(7));
    
    \count_lm_0[2]\ : CFG4
      generic map(INIT => x"D8CC")

      port map(A => un7_count_NE_i, B => count_0_sqmuxa, C => 
        count_s(2), D => state_Z(0), Y => count_lm(2));
    
    \count[24]\ : SLE
      port map(D => count_lm(24), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(24));
    
    \count[14]\ : SLE
      port map(D => count_lm(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(14));
    
    \count_lm_0[16]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(16), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(16));
    
    \tx_buffer_RNO[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(7), B => tx_buffer_Z(6), C => 
        state_Z(0), Y => N_213);
    
    \rx_data[9]\ : SLE
      port map(D => rx_buffer_Z(9), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_50_i, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_rx_data(9));
    
    \count[30]\ : SLE
      port map(D => count_lm(30), CLK => sb_sb_0_FIC_0_CLK, EN
         => N_49_i, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, SD
         => \GND\, LAT => \GND\, Q => count_Z(30));
    
    rx_data_0_sqmuxa_i_0_o3 : CFG2
      generic map(INIT => x"7")

      port map(A => un7_count_NE_i, B => state_Z(0), Y => N_320);
    
    \tx_buffer_RNO[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(3), B => tx_buffer_Z(2), C => 
        state_Z(0), Y => N_217);
    
    mosi_cl_RNO : CFG4
      generic map(INIT => x"003A")

      port map(A => \mosi_cl_0\, B => un10_count_i, C => 
        un7_count_NE_i, D => mosi_cl_4_i_0_1_Z, Y => N_25_i);
    
    assert_data : SLE
      port map(D => N_186_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        debug_led_net_0, ALn => \VCC\, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => assert_data_Z);
    
    \tx_buffer_RNO[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => spi_tx_data(11), B => tx_buffer_Z(10), C => 
        state_Z(0), Y => N_209);
    
    \count_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(11), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(10), S => count_s(11), Y => 
        count_cry_Y(11), FCO => count_cry_Z(11));
    
    \count_lm_0[20]\ : CFG3
      generic map(INIT => x"08")

      port map(A => count_s(20), B => state_Z(0), C => 
        un7_count_NE_i, Y => count_lm(20));
    
    \count_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(1), C => \GND\, D => 
        \GND\, FCI => count_s_832_FCO, S => count_s(1), Y => 
        count_cry_Y(1), FCO => count_cry_Z(1));
    
    \count_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => count_Z(9), C => \GND\, D => 
        \GND\, FCI => count_cry_Z(8), S => count_s(9), Y => 
        count_cry_Y(9), FCO => count_cry_Z(9));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity STAMP is

    port( sb_sb_0_STAMP_PADDR   : in    std_logic_vector(11 downto 2);
          STAMP_0_data_frame    : out   std_logic_vector(63 downto 0);
          sb_sb_0_STAMP_PRDATA  : out   std_logic_vector(31 downto 0);
          dataReady_0           : out   std_logic;
          sb_sb_0_STAMP_PWDATA  : in    std_logic_vector(31 downto 0);
          stamp0_spi_miso_c     : in    std_logic;
          stamp0_spi_clock_c    : out   std_logic;
          mosi_1_0              : out   std_logic;
          mosi_cl_0             : out   std_logic;
          sb_sb_0_STAMP_PSELx   : in    std_logic;
          sb_sb_0_STAMP_PENABLE : in    std_logic;
          un1_APBState_1_5      : in    std_logic;
          sb_sb_0_STAMP_PWRITE  : in    std_logic;
          sb_sb_0_STAMP_PREADY  : out   std_logic;
          debug_led_net_0       : in    std_logic;
          stamp0_spi_dms1_cs_c  : out   std_logic;
          stamp0_spi_temp_cs_c  : out   std_logic;
          stamp0_spi_dms2_cs_c  : out   std_logic;
          sb_sb_0_FIC_0_CLK     : in    std_logic;
          debug_led_net_0_arst  : in    std_logic;
          stamp0_ready_dms1_c   : in    std_logic;
          stamp0_ready_temp_c   : in    std_logic;
          stamp0_ready_dms2_c   : in    std_logic
        );

end STAMP;

architecture DEF_ARCH of STAMP is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component spi_master_1_16
    port( component_state_0      : in    std_logic := 'U';
          spi_tx_data            : in    std_logic_vector(15 downto 0) := (others => 'U');
          spi_rx_data            : out   std_logic_vector(15 downto 0);
          delay_countere         : out   std_logic;
          N_176                  : in    std_logic := 'U';
          delay_counterlde_0_0_0 : in    std_logic := 'U';
          enable                 : in    std_logic := 'U';
          spi_busy               : out   std_logic;
          mosi_cl_0              : out   std_logic;
          mosi_1_0               : out   std_logic;
          debug_led_net_0        : in    std_logic := 'U';
          stamp0_spi_clock_c     : out   std_logic;
          debug_led_net_0_arst   : in    std_logic := 'U';
          stamp0_spi_miso_c      : in    std_logic := 'U';
          sb_sb_0_FIC_0_CLK      : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \STAMP_0_data_frame\ : std_logic_vector(63 downto 0);
    signal \stamp0_spi_temp_cs_c\ : std_logic;
    signal component_state_Z : std_logic_vector(5 downto 0);
    signal async_prescaler_count_Z : 
        std_logic_vector(11 downto 0);
    signal async_prescaler_count_5_Z : 
        std_logic_vector(11 downto 0);
    signal config_Z : std_logic_vector(31 downto 3);
    signal config_RNO_0_Z : std_logic_vector(31 to 31);
    signal async_state_Z : std_logic_vector(1 downto 0);
    signal async_state_17 : std_logic_vector(1 to 1);
    signal spi_tx_data_Z : std_logic_vector(15 downto 0);
    signal spi_request_for_Z : std_logic_vector(1 downto 0);
    signal dummy_Z : std_logic_vector(31 downto 0);
    signal spi_rx_data : std_logic_vector(15 downto 0);
    signal un1_spi_rx_data_Z : std_logic_vector(14 downto 6);
    signal component_state_ns : std_logic_vector(3 downto 0);
    signal delay_counter_Z : std_logic_vector(27 downto 0);
    signal delay_counter_lm : std_logic_vector(27 downto 0);
    signal status_async_cycles_lm : std_logic_vector(5 downto 0);
    signal delay_counter_cry_Z : std_logic_vector(26 downto 0);
    signal delay_counter_cry_S : std_logic_vector(0 to 0);
    signal delay_counter_cry_Y : std_logic_vector(26 downto 0);
    signal delay_counter_s : std_logic_vector(26 downto 1);
    signal delay_counter_s_FCO : std_logic_vector(27 to 27);
    signal delay_counter_s_Z : std_logic_vector(27 to 27);
    signal delay_counter_s_Y : std_logic_vector(27 to 27);
    signal status_async_cycles_cry_Z : 
        std_logic_vector(4 downto 1);
    signal status_async_cycles_s : std_logic_vector(4 downto 1);
    signal status_async_cycles_cry_Y : 
        std_logic_vector(4 downto 1);
    signal status_async_cycles_s_FCO : std_logic_vector(5 to 5);
    signal status_async_cycles_s_Z : std_logic_vector(5 to 5);
    signal status_async_cycles_s_Y : std_logic_vector(5 to 5);
    signal un1_spi_rx_data_2_1_1_Z : 
        std_logic_vector(2 downto 0);
    signal component_state_ns_0_a3_0_0_Z : 
        std_logic_vector(0 to 0);
    signal async_state_17_iv_0_0_a3_0_1_Z : 
        std_logic_vector(1 to 1);
    signal component_state_ns_0_0_0_0_Z : 
        std_logic_vector(1 to 1);
    signal component_state_ns_0_0_0_a3_2_Z : 
        std_logic_vector(2 to 2);
    signal async_state_17_iv_0_0_0_Z : std_logic_vector(1 to 1);
    signal component_state_ns_0_0_Z : std_logic_vector(0 to 0);
    signal component_state_ns_0_0_0_a3_1_0_Z : 
        std_logic_vector(1 to 1);
    signal component_state_ns_0_1_Z : std_logic_vector(0 to 0);
    signal stamp0_ready_dms2_c_i, stamp0_ready_temp_c_i, 
        stamp0_ready_dms1_c_i, 
        un1_presetn_inv_i_a3_0_a2_0_RNINN9L1_Z, N_1454_i, N_103_i, 
        \VCC\, un5_async_prescaler_count_cry_9_S, \GND\, 
        un5_async_prescaler_count_cry_10_S, config_143, N_266_i, 
        N_33_i, un5_async_prescaler_count_cry_1_S, 
        un5_async_prescaler_count_cry_3_S, 
        un5_async_prescaler_count_cry_4_S, 
        un5_async_prescaler_count_cry_5_S, N_414_i, 
        un1_presetn_inv_2_i, N_413_i, N_570_i, 
        un1_presetn_inv_4_i, N_428_i, N_427_i, N_426_i, N_425_i, 
        N_424_i, N_423_i, N_422_i, N_421_i, N_420_i, N_419_i, 
        N_418_i, N_417_i, N_416_i, N_415_i, 
        un1_request_resync_0_sqmuxa_1_0_0_Z, N_569_i, 
        measurement_dms1_0_sqmuxa_1_Z, 
        measurement_dms2_1_sqmuxa_Z, measurement_temp_1_sqmuxa_Z, 
        un1_presetn_inv_i_a3_0_a3_Z, N_698, N_700, N_685, N_686, 
        N_687, N_688, N_689, N_690, drdy_flank_detected_temp_Z, 
        drdy_flank_detected_temp_1_sqmuxa_2_i_0_0_Z, 
        drdy_flank_detected_dms2_Z, N_21, 
        drdy_flank_detected_dms1_Z, N_23, enable, N_898, 
        un1_component_state_9_i, new_avail_0_sqmuxa_1_Z, 
        un1_new_avail_1_sqmuxa_3_i_0_0_Z, 
        request_resync_1_sqmuxa_1, N_40, 
        status_temp_overwrittenVal_9_Z, 
        un1_new_avail_0_sqmuxa_2_0_0_Z, 
        drdy_flank_detected_temp_1_sqmuxa_1, N_268_i, 
        un1_new_avail_0_sqmuxa_3_0_0_Z, 
        drdy_flank_detected_dms2_1_sqmuxa_1, N_270_i, 
        un1_drdy_flank_detected_dms1_0_sqmuxa_1_0_0_Z, 
        drdy_flank_detected_dms1_0_sqmuxa_1_Z, apb_is_reset_Z, 
        N_178_i, apb_is_atomic_Z, N_28, N_151_i, 
        spi_dms2_cs_13_iv_i_Z, N_162, spi_temp_cs_ldmx_Z, 
        N_165_tz, spi_dms1_cs_14_iv_i_Z, N_167, 
        apb_spi_finished_Z, un1_apb_spi_finished_1_f0_Z, 
        PREADY_0_sqmuxa_2, un1_PREADY_0_sqmuxa_3_0_0_Z, N_675, 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, N_676, N_677, N_678, 
        N_679, N_680, N_681, N_682, N_683, N_668, N_669, N_670, 
        N_671, N_672, N_673, N_674, delay_countere, 
        status_async_cyclese, un45_async_state_cry_0_Z, 
        un45_async_state_cry_0_S, un45_async_state_cry_0_Y, 
        un45_async_state_cry_1_Z, un45_async_state_cry_1_S, 
        un45_async_state_cry_1_Y, un45_async_state_cry_2_Z, 
        un45_async_state_cry_2_S, un45_async_state_cry_2_Y, 
        un45_async_state_cry_3_Z, un45_async_state_cry_3_S, 
        un45_async_state_cry_3_Y, un45_async_state_cry_4_Z, 
        un45_async_state_cry_4_S, un45_async_state_cry_4_Y, 
        un45_async_state_cry_5_Z, un45_async_state_cry_5_S, 
        un45_async_state_cry_5_Y, status_async_cycles_s_831_FCO, 
        status_async_cycles_s_831_S, status_async_cycles_s_831_Y, 
        un5_async_prescaler_count_s_1_837_FCO, 
        un5_async_prescaler_count_s_1_837_S, 
        un5_async_prescaler_count_s_1_837_Y, 
        un5_async_prescaler_count_cry_1_Z, 
        un5_async_prescaler_count_cry_1_Y, 
        un5_async_prescaler_count_cry_2_Z, 
        un5_async_prescaler_count_cry_2_S, 
        un5_async_prescaler_count_cry_2_Y, 
        un5_async_prescaler_count_cry_3_Z, 
        un5_async_prescaler_count_cry_3_Y, 
        un5_async_prescaler_count_cry_4_Z, 
        un5_async_prescaler_count_cry_4_Y, 
        un5_async_prescaler_count_cry_5_Z, 
        un5_async_prescaler_count_cry_5_Y, 
        un5_async_prescaler_count_cry_6_Z, 
        un5_async_prescaler_count_cry_6_S, 
        un5_async_prescaler_count_cry_6_Y, 
        un5_async_prescaler_count_cry_7_Z, 
        un5_async_prescaler_count_cry_7_S, 
        un5_async_prescaler_count_cry_7_Y, 
        un5_async_prescaler_count_cry_8_Z, 
        un5_async_prescaler_count_cry_8_S, 
        un5_async_prescaler_count_cry_8_Y, 
        un5_async_prescaler_count_cry_9_Z, 
        un5_async_prescaler_count_cry_9_Y, 
        un5_async_prescaler_count_s_11_FCO, 
        un5_async_prescaler_count_s_11_S, 
        un5_async_prescaler_count_s_11_Y, 
        un5_async_prescaler_count_cry_10_Z, 
        un5_async_prescaler_count_cry_10_Y, next_state_0_sqmuxa_Z, 
        PRDATA_684_1_Z, un1_presetn_inv_i_a3_0_a2_0_sx_Z, N_486, 
        apb_spi_finished_0_sqmuxa_1, 
        un1_presetn_inv_i_a3_0_a2_0_x_Z, N_496, 
        un1_presetn_inv_i_a3_0_a2_0_1_0_Z, 
        un1_request_resync_0_sqmuxa_1_0_0_1_Z, N_493, 
        un1_spi_rx_data_sn_N_5, N_652, N_653, N_654, 
        drdy_flank_detected_dms2_1_sqmuxa_1_0_a4_0_a3_0_Z, 
        new_avail_0_sqmuxa_1_1_Z, spi_dms2_cs_1_sqmuxa_0_Z, 
        apb_spi_finished_1_sqmuxa_0, N_378, 
        spi_dms2_cs_0_sqmuxa_Z, N_280, spi_N_5_mux_i, N_279, 
        PREADY_0_sqmuxa, N_353_i, un3_spi_busy, N_282, N_543, 
        N_594, N_593, N_592, N_591, N_601, N_614, N_616, N_595, 
        N_596, N_597, N_599, N_629, N_630, N_631, N_633, N_590, 
        N_610, N_624, N_644, N_598, N_647, N_613, N_107, N_643, 
        N_637, N_623, N_609, N_603, N_589, N_636, N_602, N_649, 
        N_615, N_588, N_600, N_622, N_634, N_635, N_604, N_605, 
        N_606, N_607, N_608, N_611, N_612, N_638, N_639, N_640, 
        N_641, N_642, N_645, N_646, un1_component_state_9_1_Z, 
        un1_component_state_9_2_0_a3_0_0, spi_busy, 
        delay_counterlde_0_0_a3_2, un27_paddr_0_0_0_1_Z, 
        N_519_i_0_a2_20, N_519_i_0_a2_19, N_519_i_0_a2_18, 
        N_519_i_0_a2_17, N_519_i_0_a2_16, N_519_i_0_a2_15, 
        N_519_i_0_a2_14, un1_async_prescaler_countlt8, N_318, 
        apb_spi_finished_1_sqmuxa_Z, un14_delay_counter_Z, 
        un15_delay_counter_Z, N_47_i_Z, next_state_1_sqmuxa, 
        N_277, N_498, spi_request_for_2_sqmuxa_Z, 
        spi_temp_cs_13_iv, spi_dms2_cs_1_sqmuxa_1_Z, N_332_i, 
        N_628, N_627, N_626, N_625, N_648, N_650, N_632, 
        un27_paddr_i_0, un1_async_prescaler_countlt10, N_662, 
        N_663, N_664, N_666, N_657, N_656, N_655, N_667, 
        spi_dms1_cs_0_sqmuxa_3_Z, spi_temp_cs_0_sqmuxa_Z, 
        N_519_i_0_a2_25, N_319, N_487, N_661, N_660, N_659, N_658, 
        N_665, un1_async_state_0_sqmuxa_i, N_331, N_309, 
        un1_async_prescaler_count, 
        status_async_cycles_2_sqmuxa_i_4, N_176, 
        status_async_cycles_1_sqmuxa_1_i_0_0_0, 
        un1_component_state_13_0_i_a3_0_1_0_Z, N_386, N_381, 
        measurement_dms1_0_sqmuxa_Z, 
        status_async_cycles_3_sqmuxa_Z, 
        status_async_cycles_2_sqmuxa_Z, N_392, 
        spi_tx_data_0_sqmuxa_Z, spi_enable_1_sqmuxa_1_Z, 
        status_async_cycles_1_sqmuxa, un1_component_state_9_3_Z, 
        un1_component_state_17_0_i_a3_0_Z, delay_counterlde_0_0_0, 
        un1_component_state_14_0_i_a3_0_s_0_Z, N_499, N_275, N_10, 
        N_9, N_8, N_7, N_6, N_5 : std_logic;

    for all : spi_master_1_16
	Use entity work.spi_master_1_16(DEF_ARCH);
begin 

    STAMP_0_data_frame(63) <= \STAMP_0_data_frame\(63);
    STAMP_0_data_frame(62) <= \STAMP_0_data_frame\(62);
    STAMP_0_data_frame(61) <= \STAMP_0_data_frame\(61);
    STAMP_0_data_frame(60) <= \STAMP_0_data_frame\(60);
    STAMP_0_data_frame(59) <= \STAMP_0_data_frame\(59);
    STAMP_0_data_frame(58) <= \STAMP_0_data_frame\(58);
    STAMP_0_data_frame(57) <= \STAMP_0_data_frame\(57);
    STAMP_0_data_frame(56) <= \STAMP_0_data_frame\(56);
    STAMP_0_data_frame(55) <= \STAMP_0_data_frame\(55);
    STAMP_0_data_frame(54) <= \STAMP_0_data_frame\(54);
    STAMP_0_data_frame(53) <= \STAMP_0_data_frame\(53);
    STAMP_0_data_frame(52) <= \STAMP_0_data_frame\(52);
    STAMP_0_data_frame(51) <= \STAMP_0_data_frame\(51);
    STAMP_0_data_frame(50) <= \STAMP_0_data_frame\(50);
    STAMP_0_data_frame(49) <= \STAMP_0_data_frame\(49);
    STAMP_0_data_frame(48) <= \STAMP_0_data_frame\(48);
    STAMP_0_data_frame(47) <= \STAMP_0_data_frame\(47);
    STAMP_0_data_frame(46) <= \STAMP_0_data_frame\(46);
    STAMP_0_data_frame(45) <= \STAMP_0_data_frame\(45);
    STAMP_0_data_frame(44) <= \STAMP_0_data_frame\(44);
    STAMP_0_data_frame(43) <= \STAMP_0_data_frame\(43);
    STAMP_0_data_frame(42) <= \STAMP_0_data_frame\(42);
    STAMP_0_data_frame(41) <= \STAMP_0_data_frame\(41);
    STAMP_0_data_frame(40) <= \STAMP_0_data_frame\(40);
    STAMP_0_data_frame(39) <= \STAMP_0_data_frame\(39);
    STAMP_0_data_frame(38) <= \STAMP_0_data_frame\(38);
    STAMP_0_data_frame(37) <= \STAMP_0_data_frame\(37);
    STAMP_0_data_frame(36) <= \STAMP_0_data_frame\(36);
    STAMP_0_data_frame(35) <= \STAMP_0_data_frame\(35);
    STAMP_0_data_frame(34) <= \STAMP_0_data_frame\(34);
    STAMP_0_data_frame(33) <= \STAMP_0_data_frame\(33);
    STAMP_0_data_frame(32) <= \STAMP_0_data_frame\(32);
    STAMP_0_data_frame(31) <= \STAMP_0_data_frame\(31);
    STAMP_0_data_frame(30) <= \STAMP_0_data_frame\(30);
    STAMP_0_data_frame(29) <= \STAMP_0_data_frame\(29);
    STAMP_0_data_frame(28) <= \STAMP_0_data_frame\(28);
    STAMP_0_data_frame(27) <= \STAMP_0_data_frame\(27);
    STAMP_0_data_frame(26) <= \STAMP_0_data_frame\(26);
    STAMP_0_data_frame(25) <= \STAMP_0_data_frame\(25);
    STAMP_0_data_frame(24) <= \STAMP_0_data_frame\(24);
    STAMP_0_data_frame(23) <= \STAMP_0_data_frame\(23);
    STAMP_0_data_frame(22) <= \STAMP_0_data_frame\(22);
    STAMP_0_data_frame(21) <= \STAMP_0_data_frame\(21);
    STAMP_0_data_frame(20) <= \STAMP_0_data_frame\(20);
    STAMP_0_data_frame(19) <= \STAMP_0_data_frame\(19);
    STAMP_0_data_frame(18) <= \STAMP_0_data_frame\(18);
    STAMP_0_data_frame(17) <= \STAMP_0_data_frame\(17);
    STAMP_0_data_frame(16) <= \STAMP_0_data_frame\(16);
    STAMP_0_data_frame(15) <= \STAMP_0_data_frame\(15);
    STAMP_0_data_frame(14) <= \STAMP_0_data_frame\(14);
    STAMP_0_data_frame(13) <= \STAMP_0_data_frame\(13);
    STAMP_0_data_frame(12) <= \STAMP_0_data_frame\(12);
    STAMP_0_data_frame(11) <= \STAMP_0_data_frame\(11);
    STAMP_0_data_frame(10) <= \STAMP_0_data_frame\(10);
    STAMP_0_data_frame(9) <= \STAMP_0_data_frame\(9);
    STAMP_0_data_frame(8) <= \STAMP_0_data_frame\(8);
    STAMP_0_data_frame(7) <= \STAMP_0_data_frame\(7);
    STAMP_0_data_frame(6) <= \STAMP_0_data_frame\(6);
    STAMP_0_data_frame(5) <= \STAMP_0_data_frame\(5);
    STAMP_0_data_frame(4) <= \STAMP_0_data_frame\(4);
    STAMP_0_data_frame(3) <= \STAMP_0_data_frame\(3);
    STAMP_0_data_frame(2) <= \STAMP_0_data_frame\(2);
    STAMP_0_data_frame(1) <= \STAMP_0_data_frame\(1);
    STAMP_0_data_frame(0) <= \STAMP_0_data_frame\(0);
    stamp0_spi_temp_cs_c <= \stamp0_spi_temp_cs_c\;

    \component_state_RNIS3IV[2]\ : CFG4
      generic map(INIT => x"0002")

      port map(A => spi_busy, B => component_state_Z(0), C => 
        component_state_Z(4), D => component_state_Z(2), Y => 
        delay_counterlde_0_0_a3_2);
    
    \delay_counter_cry[10]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(10), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(9), S => 
        delay_counter_s(10), Y => delay_counter_cry_Y(10), FCO
         => delay_counter_cry_Z(10));
    
    \measurement_temp[5]\ : SLE
      port map(D => spi_rx_data(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(21));
    
    drdy_flank_detected_temp_1_sqmuxa_1_0_a4_0_a3 : CFG3
      generic map(INIT => x"08")

      port map(A => spi_request_for_Z(1), B => 
        apb_spi_finished_0_sqmuxa_1, C => spi_request_for_Z(0), Y
         => drdy_flank_detected_temp_1_sqmuxa_1);
    
    \dummy[30]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(30));
    
    \dummy[1]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(1));
    
    \un1_spi_rx_data_0[14]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(14), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(14), Y => N_599);
    
    \async_state_17_iv_0_0_a2_RNI121S1[1]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => component_state_Z(0), B => N_282, C => 
        status_async_cycles_1_sqmuxa_1_i_0_0_0, D => N_499, Y => 
        status_async_cyclese);
    
    \delay_counter_lm_0[17]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(17), Y => 
        delay_counter_lm(17));
    
    \async_prescaler_count_5[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => un1_async_prescaler_count, B => 
        async_prescaler_count_Z(0), Y => 
        async_prescaler_count_5_Z(0));
    
    \measurement_dms1[15]\ : SLE
      port map(D => spi_rx_data(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(63));
    
    un3_spi_busy_0_a3 : CFG2
      generic map(INIT => x"1")

      port map(A => spi_request_for_Z(1), B => 
        spi_request_for_Z(0), Y => un3_spi_busy);
    
    un45_async_state_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => config_Z(24), B => \STAMP_0_data_frame\(3), C
         => \GND\, D => \GND\, FCI => \GND\, S => 
        un45_async_state_cry_0_S, Y => un45_async_state_cry_0_Y, 
        FCO => un45_async_state_cry_0_Z);
    
    new_avail_0_sqmuxa_1_1 : CFG2
      generic map(INIT => x"8")

      port map(A => component_state_Z(5), B => config_Z(30), Y
         => new_avail_0_sqmuxa_1_1_Z);
    
    \measurement_dms1[12]\ : SLE
      port map(D => spi_rx_data(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(60));
    
    \spi_request_for[0]\ : SLE
      port map(D => N_569_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_4_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_request_for_Z(0));
    
    \async_prescaler_count_5[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => un1_async_prescaler_count, B => 
        un5_async_prescaler_count_cry_7_S, Y => 
        async_prescaler_count_5_Z(7));
    
    new_avail_0_sqmuxa_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => \STAMP_0_data_frame\(15), B => 
        \STAMP_0_data_frame\(14), C => new_avail_0_sqmuxa_1_1_Z, 
        D => N_309, Y => new_avail_0_sqmuxa_1_Z);
    
    \status_async_cycles_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => \STAMP_0_data_frame\(6), C => 
        \GND\, D => \GND\, FCI => status_async_cycles_cry_Z(2), S
         => status_async_cycles_s(3), Y => 
        status_async_cycles_cry_Y(3), FCO => 
        status_async_cycles_cry_Z(3));
    
    spi_enable_RNO : CFG3
      generic map(INIT => x"EC")

      port map(A => spi_tx_data_0_sqmuxa_Z, B => 
        component_state_Z(3), C => un14_delay_counter_Z, Y => 
        N_898);
    
    \component_state_ns_0_0_0_a3_1_0[1]\ : CFG3
      generic map(INIT => x"40")

      port map(A => next_state_0_sqmuxa_Z, B => N_309, C => 
        component_state_Z(5), Y => 
        component_state_ns_0_0_0_a3_1_0_Z(1));
    
    \measurement_dms2[7]\ : SLE
      port map(D => spi_rx_data(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(39));
    
    \un1_spi_rx_data_0[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(7), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(7), Y => N_592);
    
    \config[13]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(13));
    
    \spi_tx_data_RNO[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(7), B => 
        component_state_Z(5), Y => N_421_i);
    
    \delay_counter[25]\ : SLE
      port map(D => delay_counter_lm(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(25));
    
    \dummy[27]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(27));
    
    \dummy[12]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(12));
    
    spi_dms1_cs_14_iv_i : CFG3
      generic map(INIT => x"13")

      port map(A => component_state_Z(3), B => 
        spi_dms1_cs_0_sqmuxa_3_Z, C => sb_sb_0_STAMP_PADDR(4), Y
         => spi_dms1_cs_14_iv_i_Z);
    
    \un1_spi_rx_data_1[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(37), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(5), Y => N_624);
    
    \un1_spi_rx_data_0[13]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(13), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(13), Y => N_598);
    
    un5_async_prescaler_count_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(7), C => 
        \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_6_Z, S => 
        un5_async_prescaler_count_cry_7_S, Y => 
        un5_async_prescaler_count_cry_7_Y, FCO => 
        un5_async_prescaler_count_cry_7_Z);
    
    \un1_spi_rx_data_0[16]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(16), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(16), Y => N_601);
    
    \component_state_ns_i_a3_i_0_a3_0[4]\ : CFG3
      generic map(INIT => x"40")

      port map(A => apb_spi_finished_Z, B => component_state_Z(3), 
        C => N_47_i_Z, Y => next_state_1_sqmuxa);
    
    \PRDATA[26]\ : SLE
      port map(D => N_678, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(26));
    
    measurement_dms1_0_sqmuxa_1 : CFG2
      generic map(INIT => x"8")

      port map(A => measurement_dms1_0_sqmuxa_Z, B => 
        un3_spi_busy, Y => measurement_dms1_0_sqmuxa_1_Z);
    
    \async_prescaler_count[9]\ : SLE
      port map(D => un5_async_prescaler_count_cry_9_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(9));
    
    \status_async_cycles_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => \STAMP_0_data_frame\(7), C => 
        \GND\, D => \GND\, FCI => status_async_cycles_cry_Z(3), S
         => status_async_cycles_s(4), Y => 
        status_async_cycles_cry_Y(4), FCO => 
        status_async_cycles_cry_Z(4));
    
    \spi_tx_data_RNO[15]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(15), B => 
        component_state_Z(5), Y => N_413_i);
    
    measurement_dms2_1_sqmuxa : CFG3
      generic map(INIT => x"40")

      port map(A => spi_request_for_Z(1), B => 
        measurement_dms1_0_sqmuxa_Z, C => spi_request_for_Z(0), Y
         => measurement_dms2_1_sqmuxa_Z);
    
    \spi_tx_data_RNO[11]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(11), B => 
        component_state_Z(5), Y => N_417_i);
    
    un5_async_prescaler_count_s_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(11), C
         => \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_10_Z, S => 
        un5_async_prescaler_count_s_11_S, Y => 
        un5_async_prescaler_count_s_11_Y, FCO => 
        un5_async_prescaler_count_s_11_FCO);
    
    \un1_spi_rx_data_0[24]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame\(24), B => config_Z(24), 
        C => sb_sb_0_STAMP_PADDR(8), Y => N_609);
    
    status_dms2_overwrittenVal_RNO : CFG3
      generic map(INIT => x"04")

      port map(A => N_498, B => \STAMP_0_data_frame\(14), C => 
        N_493, Y => N_268_i);
    
    \delay_counter_RNI6DFR[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => delay_counter_Z(3), B => delay_counter_Z(2), 
        C => delay_counter_Z(1), D => delay_counter_Z(0), Y => 
        N_519_i_0_a2_18);
    
    \delay_counter_lm_0[10]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(10), Y => 
        delay_counter_lm(10));
    
    \measurement_temp[4]\ : SLE
      port map(D => spi_rx_data(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(20));
    
    \async_state[1]\ : SLE
      port map(D => async_state_17(1), CLK => sb_sb_0_FIC_0_CLK, 
        EN => \VCC\, ALn => debug_led_net_0_arst, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        async_state_Z(1));
    
    apb_spi_finished : SLE
      port map(D => un1_apb_spi_finished_1_f0_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => debug_led_net_0, ALn => \VCC\, 
        ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q
         => apb_spi_finished_Z);
    
    \delay_counter[3]\ : SLE
      port map(D => delay_counter_lm(3), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(3));
    
    \async_prescaler_count[11]\ : SLE
      port map(D => async_prescaler_count_5_Z(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(11));
    
    \delay_counter[1]\ : SLE
      port map(D => delay_counter_lm(1), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(1));
    
    \spi_tx_data[15]\ : SLE
      port map(D => N_413_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(15));
    
    \status_async_cycles_lm_0[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => status_async_cycles_3_sqmuxa_Z, B => 
        status_async_cycles_s(2), C => 
        status_async_cycles_1_sqmuxa, Y => 
        status_async_cycles_lm(2));
    
    \un1_spi_rx_data_0[23]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(23), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(23), Y => N_608);
    
    \un1_spi_rx_data_0[26]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame\(26), B => config_Z(26), 
        C => sb_sb_0_STAMP_PADDR(8), Y => N_611);
    
    status_async_cycles_2_sqmuxa : CFG3
      generic map(INIT => x"80")

      port map(A => status_async_cycles_2_sqmuxa_i_4, B => 
        un3_spi_busy, C => N_309, Y => 
        status_async_cycles_2_sqmuxa_Z);
    
    \un1_spi_rx_data_2[30]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_649, B => N_615, C => N_107, Y => N_682);
    
    un5_async_prescaler_count_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(4), C => 
        \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_3_Z, S => 
        un5_async_prescaler_count_cry_4_S, Y => 
        un5_async_prescaler_count_cry_4_Y, FCO => 
        un5_async_prescaler_count_cry_4_Z);
    
    un1_new_avail_0_sqmuxa_2_0_0 : CFG3
      generic map(INIT => x"FE")

      port map(A => N_498, B => N_493, C => 
        drdy_flank_detected_temp_1_sqmuxa_1, Y => 
        un1_new_avail_0_sqmuxa_2_0_0_Z);
    
    \spi_tx_data_RNO[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(0), B => 
        component_state_Z(5), Y => N_428_i);
    
    \dummy[25]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(25));
    
    \measurement_dms2[1]\ : SLE
      port map(D => spi_rx_data(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(33));
    
    un1_request_resync_0_sqmuxa_1_0_0 : CFG4
      generic map(INIT => x"F4F0")

      port map(A => un1_request_resync_0_sqmuxa_1_0_0_1_Z, B => 
        N_486, C => N_493, D => sb_sb_0_STAMP_PADDR(8), Y => 
        un1_request_resync_0_sqmuxa_1_0_0_Z);
    
    \component_state_ns_0_0_0[1]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => component_state_ns_0_0_0_0_Z(1), B => 
        component_state_ns_0_0_0_a3_1_0_Z(1), C => 
        sb_sb_0_STAMP_PSELx, Y => component_state_ns(1));
    
    \delay_counter_lm_0[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_332_i, B => N_176, C => delay_counter_s(1), 
        Y => delay_counter_lm(1));
    
    \un1_spi_rx_data_2[18]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_637, B => N_603, C => N_107, Y => N_670);
    
    \delay_counter_cry[21]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(21), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(20), S => 
        delay_counter_s(21), Y => delay_counter_cry_Y(21), FCO
         => delay_counter_cry_Z(21));
    
    \measurement_temp[10]\ : SLE
      port map(D => spi_rx_data(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(26));
    
    un1_async_state_0_sqmuxa_0_0_0_a2 : CFG3
      generic map(INIT => x"20")

      port map(A => component_state_Z(2), B => 
        sb_sb_0_STAMP_PENABLE, C => apb_is_reset_Z, Y => N_498);
    
    \component_state[3]\ : SLE
      port map(D => component_state_ns(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => component_state_Z(3));
    
    \spi_tx_data[13]\ : SLE
      port map(D => N_415_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(13));
    
    spi : spi_master_1_16
      port map(component_state_0 => component_state_Z(5), 
        spi_tx_data(15) => spi_tx_data_Z(15), spi_tx_data(14) => 
        spi_tx_data_Z(14), spi_tx_data(13) => spi_tx_data_Z(13), 
        spi_tx_data(12) => spi_tx_data_Z(12), spi_tx_data(11) => 
        spi_tx_data_Z(11), spi_tx_data(10) => spi_tx_data_Z(10), 
        spi_tx_data(9) => spi_tx_data_Z(9), spi_tx_data(8) => 
        spi_tx_data_Z(8), spi_tx_data(7) => spi_tx_data_Z(7), 
        spi_tx_data(6) => spi_tx_data_Z(6), spi_tx_data(5) => 
        spi_tx_data_Z(5), spi_tx_data(4) => spi_tx_data_Z(4), 
        spi_tx_data(3) => spi_tx_data_Z(3), spi_tx_data(2) => 
        spi_tx_data_Z(2), spi_tx_data(1) => spi_tx_data_Z(1), 
        spi_tx_data(0) => spi_tx_data_Z(0), spi_rx_data(15) => 
        spi_rx_data(15), spi_rx_data(14) => spi_rx_data(14), 
        spi_rx_data(13) => spi_rx_data(13), spi_rx_data(12) => 
        spi_rx_data(12), spi_rx_data(11) => spi_rx_data(11), 
        spi_rx_data(10) => spi_rx_data(10), spi_rx_data(9) => 
        spi_rx_data(9), spi_rx_data(8) => spi_rx_data(8), 
        spi_rx_data(7) => spi_rx_data(7), spi_rx_data(6) => 
        spi_rx_data(6), spi_rx_data(5) => spi_rx_data(5), 
        spi_rx_data(4) => spi_rx_data(4), spi_rx_data(3) => 
        spi_rx_data(3), spi_rx_data(2) => spi_rx_data(2), 
        spi_rx_data(1) => spi_rx_data(1), spi_rx_data(0) => 
        spi_rx_data(0), delay_countere => delay_countere, N_176
         => N_176, delay_counterlde_0_0_0 => 
        delay_counterlde_0_0_0, enable => enable, spi_busy => 
        spi_busy, mosi_cl_0 => mosi_cl_0, mosi_1_0 => mosi_1_0, 
        debug_led_net_0 => debug_led_net_0, stamp0_spi_clock_c
         => stamp0_spi_clock_c, debug_led_net_0_arst => 
        debug_led_net_0_arst, stamp0_spi_miso_c => 
        stamp0_spi_miso_c, sb_sb_0_FIC_0_CLK => sb_sb_0_FIC_0_CLK);
    
    PREADY : SLE
      port map(D => PREADY_0_sqmuxa_2, CLK => sb_sb_0_FIC_0_CLK, 
        EN => un1_PREADY_0_sqmuxa_3_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => sb_sb_0_STAMP_PREADY);
    
    \PRDATA[7]\ : SLE
      port map(D => un1_spi_rx_data_Z(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_presetn_inv_i_a3_0_a3_Z, ALn
         => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => sb_sb_0_STAMP_PRDATA(7));
    
    \measurement_temp[11]\ : SLE
      port map(D => spi_rx_data(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(27));
    
    \measurement_dms1[7]\ : SLE
      port map(D => spi_rx_data(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(55));
    
    \delay_counter_lm_0[16]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(16), Y => 
        delay_counter_lm(16));
    
    \component_state[1]\ : SLE
      port map(D => N_28, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => component_state_Z(1));
    
    \un1_spi_rx_data[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_653, B => un1_spi_rx_data_sn_N_5, C => 
        spi_rx_data(1), Y => N_686);
    
    \async_state_17_iv_0_0_a3_0_1[1]\ : CFG3
      generic map(INIT => x"10")

      port map(A => component_state_Z(5), B => N_318, C => 
        async_state_Z(0), Y => async_state_17_iv_0_0_a3_0_1_Z(1));
    
    \un1_spi_rx_data_2[11]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_630, B => N_596, C => N_107, Y => N_663);
    
    \PRDATA[14]\ : SLE
      port map(D => un1_spi_rx_data_Z(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_presetn_inv_i_a3_0_a3_Z, ALn
         => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => sb_sb_0_STAMP_PRDATA(14));
    
    \config[25]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(25), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(25));
    
    \dummy[7]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(7));
    
    \un1_spi_rx_data_0[9]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(9), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(9), Y => N_594);
    
    \dummy[17]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(17));
    
    \un1_spi_rx_data_1[22]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(54), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(22), Y => N_641);
    
    \config[7]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(7));
    
    \component_state[2]\ : SLE
      port map(D => component_state_ns(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => component_state_Z(2));
    
    \un1_spi_rx_data_2[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_626, B => N_107, C => N_592, Y => N_659);
    
    \measurement_temp[7]\ : SLE
      port map(D => spi_rx_data(7), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(23));
    
    \measurement_dms2[6]\ : SLE
      port map(D => spi_rx_data(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(38));
    
    \async_prescaler_count[10]\ : SLE
      port map(D => un5_async_prescaler_count_cry_10_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(10));
    
    \measurement_dms1[13]\ : SLE
      port map(D => spi_rx_data(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(61));
    
    \delay_counter[5]\ : SLE
      port map(D => delay_counter_lm(5), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(5));
    
    \spi_tx_data_RNO[9]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(9), B => 
        component_state_Z(5), Y => N_419_i);
    
    \delay_counter_cry[23]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(23), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(22), S => 
        delay_counter_s(23), Y => delay_counter_cry_Y(23), FCO
         => delay_counter_cry_Z(23));
    
    \config[3]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(3));
    
    \PRDATA[27]\ : SLE
      port map(D => N_679, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(27));
    
    \delay_counter_lm_0[18]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(18), Y => 
        delay_counter_lm(18));
    
    \measurement_dms2[5]\ : SLE
      port map(D => spi_rx_data(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(37));
    
    \config[21]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(21));
    
    \un1_spi_rx_data_2[29]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_648, B => N_614, C => N_107, Y => N_681);
    
    \measurement_dms2[10]\ : SLE
      port map(D => spi_rx_data(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(42));
    
    \status_async_cycles_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => \STAMP_0_data_frame\(4), C => 
        \GND\, D => \GND\, FCI => status_async_cycles_s_831_FCO, 
        S => status_async_cycles_s(1), Y => 
        status_async_cycles_cry_Y(1), FCO => 
        status_async_cycles_cry_Z(1));
    
    \delay_counter[15]\ : SLE
      port map(D => delay_counter_lm(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(15));
    
    \un1_spi_rx_data_2_1_1[0]\ : CFG4
      generic map(INIT => x"5553")

      port map(A => \STAMP_0_data_frame\(0), B => 
        \STAMP_0_data_frame\(32), C => sb_sb_0_STAMP_PADDR(9), D
         => sb_sb_0_STAMP_PADDR(7), Y => 
        un1_spi_rx_data_2_1_1_Z(0));
    
    \config[4]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(4));
    
    \PRDATA[28]\ : SLE
      port map(D => N_680, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(28));
    
    \un1_spi_rx_data_2[20]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_639, B => N_605, C => N_107, Y => N_672);
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    \un1_spi_rx_data_1[12]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(44), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(12), Y => N_631);
    
    \delay_counter_s[27]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => \VCC\, B => delay_counter_Z(27), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(26), S => 
        delay_counter_s_Z(27), Y => delay_counter_s_Y(27), FCO
         => delay_counter_s_FCO(27));
    
    \config_RNO_0[31]\ : CFG4
      generic map(INIT => x"CCDC")

      port map(A => sb_sb_0_STAMP_PADDR(7), B => N_378, C => 
        N_496, D => sb_sb_0_STAMP_PADDR(8), Y => 
        config_RNO_0_Z(31));
    
    \un1_spi_rx_data_1[25]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(57), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(25), Y => N_644);
    
    \spi_tx_data[11]\ : SLE
      port map(D => N_417_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(11));
    
    un27_paddr_0_0_0 : CFG4
      generic map(INIT => x"F2FF")

      port map(A => sb_sb_0_STAMP_PADDR(4), B => 
        stamp0_ready_dms1_c, C => un27_paddr_0_0_0_1_Z, D => 
        sb_sb_0_STAMP_PADDR(7), Y => un27_paddr_i_0);
    
    spi_dms2_cs_1_sqmuxa_0 : CFG2
      generic map(INIT => x"4")

      port map(A => drdy_flank_detected_dms1_Z, B => 
        drdy_flank_detected_dms2_Z, Y => spi_dms2_cs_1_sqmuxa_0_Z);
    
    \measurement_dms2[11]\ : SLE
      port map(D => spi_rx_data(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(43));
    
    \component_state_ns_0_0[0]\ : CFG4
      generic map(INIT => x"30BA")

      port map(A => N_543, B => apb_is_atomic_Z, C => 
        PREADY_0_sqmuxa, D => N_309, Y => 
        component_state_ns_0_0_Z(0));
    
    \un1_spi_rx_data[8]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_660, C => 
        spi_rx_data(8), Y => un1_spi_rx_data_Z(8));
    
    \un1_spi_rx_data_1[27]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(59), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(27), Y => N_646);
    
    \un1_spi_rx_data_2[8]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_627, B => N_107, C => N_593, Y => N_660);
    
    \delay_counter[6]\ : SLE
      port map(D => delay_counter_lm(6), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(6));
    
    \config[12]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(12));
    
    \dummy[15]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(15));
    
    drdy_flank_detected_temp_RNO : CFG1
      generic map(INIT => "01")

      port map(A => stamp0_ready_temp_c, Y => 
        stamp0_ready_temp_c_i);
    
    \delay_counter[22]\ : SLE
      port map(D => delay_counter_lm(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(22));
    
    \measurement_temp[6]\ : SLE
      port map(D => spi_rx_data(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(22));
    
    \delay_counter_cry[15]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(15), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(14), S => 
        delay_counter_s(15), Y => delay_counter_cry_Y(15), FCO
         => delay_counter_cry_Z(15));
    
    \un1_spi_rx_data_0[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(4), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(4), Y => N_589);
    
    status_async_cycles_2_sqmuxa_4 : CFG4
      generic map(INIT => x"1000")

      port map(A => async_state_Z(1), B => spi_busy, C => 
        component_state_Z(0), D => un1_async_prescaler_count, Y
         => status_async_cycles_2_sqmuxa_i_4);
    
    \delay_counter_cry[16]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(16), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(15), S => 
        delay_counter_s(16), Y => delay_counter_cry_Y(16), FCO
         => delay_counter_cry_Z(16));
    
    un1_component_state_14_0_i_a3_0_s_0 : CFG4
      generic map(INIT => x"0010")

      port map(A => spi_request_for_Z(1), B => 
        spi_request_for_Z(0), C => N_309, D => spi_busy, Y => 
        un1_component_state_14_0_i_a3_0_s_0_Z);
    
    \un1_spi_rx_data_1[15]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(47), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(15), Y => N_634);
    
    \delay_counter_lm_0[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_332_i, B => N_176, C => delay_counter_s(4), 
        Y => delay_counter_lm(4));
    
    \PRDATA[10]\ : SLE
      port map(D => un1_spi_rx_data_Z(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_presetn_inv_i_a3_0_a3_Z, ALn
         => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => sb_sb_0_STAMP_PRDATA(10));
    
    \un1_spi_rx_data_1[17]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(49), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(17), Y => N_636);
    
    \component_state_ns_0_0_0_0[1]\ : CFG4
      generic map(INIT => x"AE0C")

      port map(A => apb_is_atomic_Z, B => component_state_Z(4), C
         => sb_sb_0_STAMP_PENABLE, D => PREADY_0_sqmuxa, Y => 
        component_state_ns_0_0_0_0_Z(1));
    
    \status_async_cycles_lm_0[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => status_async_cycles_3_sqmuxa_Z, B => 
        status_async_cycles_s(1), C => 
        status_async_cycles_1_sqmuxa, Y => 
        status_async_cycles_lm(1));
    
    un1_presetn_inv_i_a3_0_o2 : CFG3
      generic map(INIT => x"9E")

      port map(A => sb_sb_0_STAMP_PADDR(8), B => 
        sb_sb_0_STAMP_PADDR(7), C => sb_sb_0_STAMP_PADDR(9), Y
         => N_319);
    
    \config[20]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(20));
    
    drdy_flank_detected_dms1_RNO : CFG1
      generic map(INIT => "01")

      port map(A => stamp0_ready_dms1_c, Y => 
        stamp0_ready_dms1_c_i);
    
    \delay_counter[21]\ : SLE
      port map(D => delay_counter_lm(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(21));
    
    new_avail : SLE
      port map(D => new_avail_0_sqmuxa_1_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_new_avail_1_sqmuxa_3_i_0_0_Z, 
        ALn => debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => dataReady_0);
    
    \config[16]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(16));
    
    \PRDATA[13]\ : SLE
      port map(D => N_698, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_Z, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_STAMP_PRDATA(13));
    
    \measurement_dms1[0]\ : SLE
      port map(D => spi_rx_data(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(48));
    
    \measurement_dms1[14]\ : SLE
      port map(D => spi_rx_data(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(62));
    
    \delay_counter_lm_0[25]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(25), Y => 
        delay_counter_lm(25));
    
    status_temp_newVal : SLE
      port map(D => drdy_flank_detected_temp_1_sqmuxa_1, CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_new_avail_0_sqmuxa_2_0_0_Z, 
        ALn => debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(13));
    
    \delay_counter_cry[14]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(14), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(13), S => 
        delay_counter_s(14), Y => delay_counter_cry_Y(14), FCO
         => delay_counter_cry_Z(14));
    
    \dummy[2]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(2));
    
    \un1_spi_rx_data_0[30]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame\(30), B => config_Z(30), 
        C => sb_sb_0_STAMP_PADDR(8), Y => N_615);
    
    \PRDATA[3]\ : SLE
      port map(D => N_688, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_Z, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_STAMP_PRDATA(3));
    
    \delay_counter_cry[12]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(12), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(11), S => 
        delay_counter_s(12), Y => delay_counter_cry_Y(12), FCO
         => delay_counter_cry_Z(12));
    
    \component_state_ns_0_0_0[3]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => PREADY_0_sqmuxa_2, B => component_state_Z(2), 
        C => sb_sb_0_STAMP_PENABLE, Y => component_state_ns(3));
    
    \PRDATA[5]\ : SLE
      port map(D => N_690, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_Z, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_STAMP_PRDATA(5));
    
    \un1_spi_rx_data[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_656, C => 
        spi_rx_data(4), Y => N_689);
    
    \un1_spi_rx_data_1[31]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame\(63), B => dummy_Z(31), C
         => sb_sb_0_STAMP_PADDR(8), D => sb_sb_0_STAMP_PADDR(9), 
        Y => N_650);
    
    un27_paddr_0_0_0_1 : CFG4
      generic map(INIT => x"7530")

      port map(A => stamp0_ready_dms2_c, B => stamp0_ready_temp_c, 
        C => sb_sb_0_STAMP_PADDR(6), D => sb_sb_0_STAMP_PADDR(5), 
        Y => un27_paddr_0_0_0_1_Z);
    
    un1_PREADY_0_sqmuxa_3_0_0 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => component_state_Z(4), B => 
        component_state_Z(5), C => PREADY_0_sqmuxa, D => 
        PREADY_0_sqmuxa_2, Y => un1_PREADY_0_sqmuxa_3_0_0_Z);
    
    \measurement_temp[8]\ : SLE
      port map(D => spi_rx_data(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(24));
    
    status_async_cycles_3_sqmuxa : CFG4
      generic map(INIT => x"0080")

      port map(A => N_309, B => status_async_cycles_2_sqmuxa_i_4, 
        C => spi_request_for_Z(0), D => spi_request_for_Z(1), Y
         => status_async_cycles_3_sqmuxa_Z);
    
    \status_async_cycles[4]\ : SLE
      port map(D => status_async_cycles_lm(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => status_async_cyclese, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(7));
    
    \spi_tx_data_RNO[14]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(14), B => 
        component_state_Z(5), Y => N_414_i);
    
    \spi_tx_data_RNO[6]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(6), B => 
        component_state_Z(5), Y => N_422_i);
    
    un1_async_prescaler_countlto5 : CFG4
      generic map(INIT => x"0001")

      port map(A => async_prescaler_count_Z(5), B => 
        async_prescaler_count_Z(4), C => 
        async_prescaler_count_Z(3), D => 
        async_prescaler_count_Z(2), Y => 
        un1_async_prescaler_countlt8);
    
    \un1_spi_rx_data_0[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(6), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(6), Y => N_591);
    
    \dummy[31]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(31), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(31));
    
    status_dms2_overwrittenVal : SLE
      port map(D => N_268_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_new_avail_0_sqmuxa_3_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(11));
    
    \component_state_RNI8I9S[1]\ : CFG4
      generic map(INIT => x"0105")

      port map(A => component_state_Z(1), B => apb_spi_finished_Z, 
        C => component_state_Z(4), D => component_state_Z(3), Y
         => un1_component_state_9_2_0_a3_0_0);
    
    un1_new_avail_0_sqmuxa_3_0_0 : CFG3
      generic map(INIT => x"FE")

      port map(A => N_498, B => N_493, C => 
        drdy_flank_detected_dms2_1_sqmuxa_1, Y => 
        un1_new_avail_0_sqmuxa_3_0_0_Z);
    
    request_resync : SLE
      port map(D => request_resync_1_sqmuxa_1, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_40, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(9));
    
    \measurement_temp[3]\ : SLE
      port map(D => spi_rx_data(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(19));
    
    \delay_counter_cry[19]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(19), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(18), S => 
        delay_counter_s(19), Y => delay_counter_cry_Y(19), FCO
         => delay_counter_cry_Z(19));
    
    \un1_spi_rx_data_2[12]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_631, B => N_597, C => N_107, Y => N_664);
    
    \spi_tx_data_RNO[12]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(12), B => 
        component_state_Z(5), Y => N_416_i);
    
    \un1_spi_rx_data_0[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(5), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(5), Y => N_590);
    
    \spi_tx_data[2]\ : SLE
      port map(D => N_426_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(2));
    
    spi_enable_1_sqmuxa_1 : CFG3
      generic map(INIT => x"13")

      port map(A => N_309, B => N_282, C => next_state_0_sqmuxa_Z, 
        Y => spi_enable_1_sqmuxa_1_Z);
    
    \measurement_dms2[9]\ : SLE
      port map(D => spi_rx_data(9), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(41));
    
    \PRDATA[15]\ : SLE
      port map(D => N_700, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_Z, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_STAMP_PRDATA(15));
    
    \async_state_RNIGA801[1]\ : CFG4
      generic map(INIT => x"03AB")

      port map(A => N_493, B => un1_async_prescaler_count, C => 
        async_state_Z(1), D => component_state_Z(0), Y => 
        status_async_cycles_1_sqmuxa_1_i_0_0_0);
    
    \measurement_dms2[3]\ : SLE
      port map(D => spi_rx_data(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(35));
    
    \spi_tx_data_RNO[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(1), B => 
        component_state_Z(5), Y => N_427_i);
    
    \async_prescaler_count[1]\ : SLE
      port map(D => un5_async_prescaler_count_cry_1_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(1));
    
    \PRDATA[6]\ : SLE
      port map(D => un1_spi_rx_data_Z(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_presetn_inv_i_a3_0_a3_Z, ALn
         => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => sb_sb_0_STAMP_PRDATA(6));
    
    \delay_counter[8]\ : SLE
      port map(D => delay_counter_lm(8), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(8));
    
    \measurement_temp[2]\ : SLE
      port map(D => spi_rx_data(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(18));
    
    \spi_tx_data_RNO[8]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(8), B => 
        component_state_Z(5), Y => N_420_i);
    
    \delay_counter_lm_0[6]\ : CFG4
      generic map(INIT => x"FCAC")

      port map(A => N_332_i, B => delay_counter_s(6), C => N_176, 
        D => apb_spi_finished_0_sqmuxa_1, Y => 
        delay_counter_lm(6));
    
    drdy_flank_detected_dms1_1_sqmuxa_1_i_0_0 : CFG3
      generic map(INIT => x"FB")

      port map(A => drdy_flank_detected_dms1_0_sqmuxa_1_Z, B => 
        stamp0_ready_dms1_c, C => N_493, Y => N_23);
    
    \config[17]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(17));
    
    \delay_counter_lm_0[21]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(21), Y => 
        delay_counter_lm(21));
    
    \delay_counter[12]\ : SLE
      port map(D => delay_counter_lm(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(12));
    
    \measurement_dms1[8]\ : SLE
      port map(D => spi_rx_data(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(56));
    
    \un1_spi_rx_data[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_654, B => un1_spi_rx_data_sn_N_5, C => 
        spi_rx_data(2), Y => N_687);
    
    \status_async_cycles_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => \STAMP_0_data_frame\(5), C => 
        \GND\, D => \GND\, FCI => status_async_cycles_cry_Z(1), S
         => status_async_cycles_s(2), Y => 
        status_async_cycles_cry_Y(2), FCO => 
        status_async_cycles_cry_Z(2));
    
    \config[18]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(18));
    
    \config[2]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(2));
    
    \async_state_17_iv_0_0_o2[1]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => component_state_Z(2), B => 
        component_state_Z(3), C => component_state_Z(1), D => 
        component_state_Z(4), Y => N_318);
    
    \measurement_dms2[15]\ : SLE
      port map(D => spi_rx_data(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(47));
    
    \dummy[6]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(6));
    
    \measurement_dms2[12]\ : SLE
      port map(D => spi_rx_data(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(44));
    
    \delay_counter[19]\ : SLE
      port map(D => delay_counter_lm(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(19));
    
    \un1_spi_rx_data_2[15]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_634, B => N_600, C => N_107, Y => N_667);
    
    \config[29]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(29));
    
    \un1_spi_rx_data_2[17]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_636, B => N_602, C => N_107, Y => N_669);
    
    \spi_tx_data[3]\ : SLE
      port map(D => N_425_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(3));
    
    \un1_spi_rx_data_2[24]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_643, B => N_609, C => N_107, Y => N_676);
    
    \un1_spi_rx_data_0[18]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(18), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(18), Y => N_603);
    
    \config[14]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(14));
    
    apb_is_reset : SLE
      port map(D => sb_sb_0_STAMP_PADDR(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_178_i, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        apb_is_reset_Z);
    
    un1_request_resync_0_sqmuxa_1_0_a2_1 : CFG4
      generic map(INIT => x"0080")

      port map(A => sb_sb_0_STAMP_PADDR(9), B => 
        sb_sb_0_STAMP_PWRITE, C => 
        un1_presetn_inv_i_a3_0_a2_0_x_Z, D => un1_APBState_1_5, Y
         => N_496);
    
    un14_delay_counter : CFG3
      generic map(INIT => x"FE")

      port map(A => drdy_flank_detected_temp_Z, B => 
        drdy_flank_detected_dms2_Z, C => 
        drdy_flank_detected_dms1_Z, Y => un14_delay_counter_Z);
    
    spi_temp_cs : SLE
      port map(D => spi_temp_cs_ldmx_Z, CLK => sb_sb_0_FIC_0_CLK, 
        EN => N_165_tz, ALn => debug_led_net_0_arst, ADn => \GND\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \stamp0_spi_temp_cs_c\);
    
    \delay_counter_lm_0[13]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(13), Y => 
        delay_counter_lm(13));
    
    \delay_counter[11]\ : SLE
      port map(D => delay_counter_lm(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(11));
    
    un45_async_state_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => config_Z(25), B => \STAMP_0_data_frame\(4), C
         => \GND\, D => \GND\, FCI => un45_async_state_cry_0_Z, S
         => un45_async_state_cry_1_S, Y => 
        un45_async_state_cry_1_Y, FCO => un45_async_state_cry_1_Z);
    
    un1_PREADY_0_sqmuxa_3_0_0_a3 : CFG4
      generic map(INIT => x"8C0C")

      port map(A => apb_spi_finished_Z, B => component_state_Z(3), 
        C => N_47_i_Z, D => un27_paddr_i_0, Y => 
        PREADY_0_sqmuxa_2);
    
    \measurement_dms1[9]\ : SLE
      port map(D => spi_rx_data(9), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(57));
    
    un5_async_prescaler_count_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(10), C
         => \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_9_Z, S => 
        un5_async_prescaler_count_cry_10_S, Y => 
        un5_async_prescaler_count_cry_10_Y, FCO => 
        un5_async_prescaler_count_cry_10_Z);
    
    \un1_spi_rx_data_2[23]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_642, B => N_608, C => N_107, Y => N_675);
    
    un1_async_prescaler_countlto8 : CFG4
      generic map(INIT => x"DFFF")

      port map(A => async_prescaler_count_Z(6), B => 
        un1_async_prescaler_countlt8, C => 
        async_prescaler_count_Z(8), D => 
        async_prescaler_count_Z(7), Y => 
        un1_async_prescaler_countlt10);
    
    \un1_spi_rx_data_0[11]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(11), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(11), Y => N_596);
    
    \PRDATA[12]\ : SLE
      port map(D => un1_spi_rx_data_Z(12), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_presetn_inv_i_a3_0_a3_Z, ALn
         => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => sb_sb_0_STAMP_PRDATA(12));
    
    measurement_temp_1_sqmuxa : CFG4
      generic map(INIT => x"0800")

      port map(A => apb_spi_finished_0_sqmuxa_1, B => 
        debug_led_net_0, C => spi_request_for_Z(0), D => 
        spi_request_for_Z(1), Y => measurement_temp_1_sqmuxa_Z);
    
    \un1_spi_rx_data_2[26]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_645, B => N_611, C => N_107, Y => N_678);
    
    un1_async_prescaler_countlto11 : CFG4
      generic map(INIT => x"0F4F")

      port map(A => async_prescaler_count_Z(9), B => 
        un1_async_prescaler_countlt10, C => 
        async_prescaler_count_Z(11), D => 
        async_prescaler_count_Z(10), Y => 
        un1_async_prescaler_count);
    
    \PRDATA[19]\ : SLE
      port map(D => N_671, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(19));
    
    \dummy[20]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(20));
    
    apb_spi_finished_1_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => apb_spi_finished_0_sqmuxa_1, B => 
        apb_spi_finished_1_sqmuxa_0, Y => 
        apb_spi_finished_1_sqmuxa_Z);
    
    \dummy[0]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(0));
    
    spi_enable : SLE
      port map(D => N_898, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_component_state_9_i, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        enable);
    
    \delay_counter_cry[1]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(1), C => \GND\, D
         => \GND\, FCI => delay_counter_cry_Z(0), S => 
        delay_counter_s(1), Y => delay_counter_cry_Y(1), FCO => 
        delay_counter_cry_Z(1));
    
    \un1_spi_rx_data_0[28]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame\(28), B => config_Z(28), 
        C => sb_sb_0_STAMP_PADDR(8), Y => N_613);
    
    status_dms1_overwrittenVal_RNO : CFG3
      generic map(INIT => x"04")

      port map(A => N_498, B => \STAMP_0_data_frame\(15), C => 
        N_493, Y => N_270_i);
    
    \config[9]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(9));
    
    spi_dms1_cs : SLE
      port map(D => spi_dms1_cs_14_iv_i_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_167, ALn => 
        debug_led_net_0_arst, ADn => \GND\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => stamp0_spi_dms1_cs_c);
    
    \delay_counter[24]\ : SLE
      port map(D => delay_counter_lm(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(24));
    
    \dummy[4]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(4), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(4));
    
    un1_component_state_17_0_i_o2_0 : CFG2
      generic map(INIT => x"D")

      port map(A => spi_dms2_cs_0_sqmuxa_Z, B => config_Z(31), Y
         => N_280);
    
    drdy_flank_detected_temp_1_sqmuxa_1_0_a4_0_a3_1 : CFG3
      generic map(INIT => x"40")

      port map(A => spi_busy, B => component_state_Z(0), C => 
        N_309, Y => apb_spi_finished_0_sqmuxa_1);
    
    \delay_counter[2]\ : SLE
      port map(D => delay_counter_lm(2), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(2));
    
    \spi_tx_data_RNO[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(2), B => 
        component_state_Z(5), Y => N_426_i);
    
    \config[31]\ : SLE
      port map(D => N_266_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        config_RNO_0_Z(31), ALn => debug_led_net_0_arst, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        config_Z(31));
    
    un1_component_state_17_0_i_o2_2 : CFG3
      generic map(INIT => x"57")

      port map(A => component_state_Z(2), B => 
        sb_sb_0_STAMP_PENABLE, C => apb_is_atomic_Z, Y => N_277);
    
    \un1_spi_rx_data_0[21]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(21), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(21), Y => N_606);
    
    \PRDATA[21]\ : SLE
      port map(D => N_673, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(21));
    
    \un1_spi_rx_data_2[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_622, B => N_588, C => N_107, Y => N_655);
    
    \component_state_ns_0_a2[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => component_state_Z(5), B => 
        component_state_Z(0), Y => N_543);
    
    apb_is_atomic : SLE
      port map(D => sb_sb_0_STAMP_PADDR(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_178_i, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        apb_is_atomic_Z);
    
    \delay_counter_cry[0]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(0), C => \GND\, D
         => \GND\, FCI => \GND\, S => delay_counter_cry_S(0), Y
         => delay_counter_cry_Y(0), FCO => delay_counter_cry_Z(0));
    
    \un1_spi_rx_data_1[29]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame\(61), B => dummy_Z(29), C
         => sb_sb_0_STAMP_PADDR(8), D => sb_sb_0_STAMP_PADDR(9), 
        Y => N_648);
    
    \un1_spi_rx_data_1[20]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(52), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(20), Y => N_639);
    
    \un1_spi_rx_data_0[8]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(8), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(8), Y => N_593);
    
    \delay_counter_RNIIFLA[12]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => delay_counter_Z(15), B => delay_counter_Z(14), 
        C => delay_counter_Z(13), D => delay_counter_Z(12), Y => 
        N_519_i_0_a2_19);
    
    \delay_counter[23]\ : SLE
      port map(D => delay_counter_lm(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(23));
    
    \PRDATA[1]\ : SLE
      port map(D => N_686, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_Z, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_STAMP_PRDATA(1));
    
    \delay_counter[20]\ : SLE
      port map(D => delay_counter_lm(20), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(20));
    
    un1_apb_spi_finished_1_f0 : CFG3
      generic map(INIT => x"54")

      port map(A => N_353_i, B => apb_spi_finished_Z, C => 
        apb_spi_finished_1_sqmuxa_Z, Y => 
        un1_apb_spi_finished_1_f0_Z);
    
    un45_async_state_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => config_Z(26), B => \STAMP_0_data_frame\(5), C
         => \GND\, D => \GND\, FCI => un45_async_state_cry_1_Z, S
         => un45_async_state_cry_2_S, Y => 
        un45_async_state_cry_2_Y, FCO => un45_async_state_cry_2_Z);
    
    \dummy[24]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(24));
    
    \delay_counter_lm_0[19]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(19), Y => 
        delay_counter_lm(19));
    
    \spi_tx_data_RNO[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(3), B => 
        component_state_Z(5), Y => N_425_i);
    
    un45_async_state_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => config_Z(29), B => \STAMP_0_data_frame\(8), C
         => \GND\, D => \GND\, FCI => un45_async_state_cry_4_Z, S
         => un45_async_state_cry_5_S, Y => 
        un45_async_state_cry_5_Y, FCO => un45_async_state_cry_5_Z);
    
    un45_async_state_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => config_Z(28), B => \STAMP_0_data_frame\(7), C
         => \GND\, D => \GND\, FCI => un45_async_state_cry_3_Z, S
         => un45_async_state_cry_4_S, Y => 
        un45_async_state_cry_4_Y, FCO => un45_async_state_cry_4_Z);
    
    \component_state_RNIFR114[0]\ : CFG3
      generic map(INIT => x"CD")

      port map(A => component_state_Z(5), B => N_309, C => 
        component_state_Z(0), Y => N_176);
    
    \un1_spi_rx_data[12]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_664, C => 
        spi_rx_data(12), Y => un1_spi_rx_data_Z(12));
    
    \spi_tx_data_RNO[13]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(13), B => 
        component_state_Z(5), Y => N_415_i);
    
    PREADY_0_sqmuxa_0_a4_0_a2 : CFG2
      generic map(INIT => x"4")

      port map(A => sb_sb_0_STAMP_PENABLE, B => 
        component_state_Z(2), Y => PREADY_0_sqmuxa);
    
    \un1_spi_rx_data_1[6]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame\(38), B => dummy_Z(6), C
         => sb_sb_0_STAMP_PADDR(8), D => sb_sb_0_STAMP_PADDR(9), 
        Y => N_625);
    
    \PRDATA[31]\ : SLE
      port map(D => N_683, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(31));
    
    \config_RNO_1[31]\ : CFG2
      generic map(INIT => x"2")

      port map(A => component_state_Z(5), B => 
        component_state_Z(3), Y => N_378);
    
    \un1_spi_rx_data_1[19]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(51), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(19), Y => N_638);
    
    \un1_spi_rx_data_1[10]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(42), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(10), Y => N_629);
    
    \measurement_dms2[13]\ : SLE
      port map(D => spi_rx_data(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(45));
    
    \component_state_RNI2G06[5]\ : CFG1
      generic map(INIT => "01")

      port map(A => component_state_Z(5), Y => N_103_i);
    
    \PRDATA[16]\ : SLE
      port map(D => N_668, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(16));
    
    \delay_counter_lm_0[22]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(22), Y => 
        delay_counter_lm(22));
    
    \delay_counter[9]\ : SLE
      port map(D => delay_counter_lm(9), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(9));
    
    \config[30]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(30), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(30));
    
    un5_async_prescaler_count_s_1_837 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(0), C => 
        \GND\, D => \GND\, FCI => \VCC\, S => 
        un5_async_prescaler_count_s_1_837_S, Y => 
        un5_async_prescaler_count_s_1_837_Y, FCO => 
        un5_async_prescaler_count_s_1_837_FCO);
    
    \async_prescaler_count[2]\ : SLE
      port map(D => async_prescaler_count_5_Z(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(2));
    
    \delay_counter_lm_0[7]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(7), Y => 
        delay_counter_lm(7));
    
    \spi_tx_data[6]\ : SLE
      port map(D => N_422_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(6));
    
    un1_component_state_17_0_i_o2_2_RNI33C72 : CFG4
      generic map(INIT => x"8A00")

      port map(A => N_277, B => N_47_i_Z, C => 
        component_state_Z(3), D => 
        un1_component_state_9_2_0_a3_0_0, Y => N_487);
    
    un15_delay_counter : CFG3
      generic map(INIT => x"02")

      port map(A => drdy_flank_detected_temp_Z, B => 
        drdy_flank_detected_dms2_Z, C => 
        drdy_flank_detected_dms1_Z, Y => un15_delay_counter_Z);
    
    un1_component_state_17_0_i : CFG4
      generic map(INIT => x"D000")

      port map(A => component_state_Z(0), B => 
        un1_component_state_17_0_i_a3_0_Z, C => N_280, D => N_487, 
        Y => N_162);
    
    \dummy[10]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(10));
    
    \config_RNIMG4L[31]\ : CFG2
      generic map(INIT => x"D")

      port map(A => component_state_Z(5), B => config_Z(31), Y
         => N_282);
    
    \config[15]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(15), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(15));
    
    \PRDATA[2]\ : SLE
      port map(D => N_687, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_Z, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_STAMP_PRDATA(2));
    
    \delay_counter_cry[11]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(11), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(10), S => 
        delay_counter_s(11), Y => delay_counter_cry_Y(11), FCO
         => delay_counter_cry_Z(11));
    
    un14_delay_counter_RNIVTTH : CFG4
      generic map(INIT => x"C888")

      port map(A => next_state_1_sqmuxa, B => debug_led_net_0, C
         => un14_delay_counter_Z, D => spi_tx_data_0_sqmuxa_Z, Y
         => un1_presetn_inv_4_i);
    
    un1_new_avail_1_sqmuxa_3_i_0_0 : CFG4
      generic map(INIT => x"FEFA")

      port map(A => N_493, B => component_state_Z(5), C => N_498, 
        D => N_309, Y => un1_new_avail_1_sqmuxa_3_i_0_0_Z);
    
    \spi_tx_data[1]\ : SLE
      port map(D => N_427_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(1));
    
    \component_state_ns_0[0]\ : CFG4
      generic map(INIT => x"CCDC")

      port map(A => sb_sb_0_STAMP_PSELx, B => 
        component_state_ns_0_1_Z(0), C => N_543, D => 
        next_state_0_sqmuxa_Z, Y => component_state_ns(0));
    
    spi_dms2_cs_1_sqmuxa_1 : CFG4
      generic map(INIT => x"8000")

      port map(A => spi_dms2_cs_1_sqmuxa_0_Z, B => N_309, C => 
        config_Z(30), D => component_state_Z(5), Y => 
        spi_dms2_cs_1_sqmuxa_1_Z);
    
    \dummy[29]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(29), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(29));
    
    \un1_spi_rx_data_2[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_624, B => N_590, C => N_107, Y => N_657);
    
    \spi_request_for_RNO[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => spi_request_for_2_sqmuxa_Z, B => 
        component_state_Z(3), Y => N_570_i);
    
    \delay_counter_lm_0[24]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(24), Y => 
        delay_counter_lm(24));
    
    \status_async_cycles[1]\ : SLE
      port map(D => status_async_cycles_lm(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => status_async_cyclese, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(4));
    
    \async_state_17_iv_0_0_o2_2[1]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => component_state_Z(5), B => N_318, C => 
        async_state_Z(0), D => component_state_Z(0), Y => N_331);
    
    \delay_counter_lm_0[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(8), Y => 
        delay_counter_lm(8));
    
    un1_component_state_13_0_i_a3_0_1_0 : CFG4
      generic map(INIT => x"0020")

      port map(A => spi_request_for_Z(1), B => 
        spi_request_for_Z(0), C => N_309, D => spi_busy, Y => 
        un1_component_state_13_0_i_a3_0_1_0_Z);
    
    \delay_counter[26]\ : SLE
      port map(D => delay_counter_lm(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(26));
    
    \config[11]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(11));
    
    \delay_counter_cry[6]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(6), C => \GND\, D
         => \GND\, FCI => delay_counter_cry_Z(5), S => 
        delay_counter_s(6), Y => delay_counter_cry_Y(6), FCO => 
        delay_counter_cry_Z(6));
    
    \un1_spi_rx_data_2[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_625, B => N_107, C => N_591, Y => N_658);
    
    config_143_0_0_a4_0_a3 : CFG4
      generic map(INIT => x"0100")

      port map(A => component_state_Z(5), B => 
        sb_sb_0_STAMP_PADDR(7), C => sb_sb_0_STAMP_PADDR(8), D
         => N_496, Y => config_143);
    
    \un1_spi_rx_data[14]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_666, C => 
        spi_rx_data(14), Y => un1_spi_rx_data_Z(14));
    
    \status_async_cycles[5]\ : SLE
      port map(D => status_async_cycles_lm(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => status_async_cyclese, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(8));
    
    un5_async_prescaler_count_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(9), C => 
        \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_8_Z, S => 
        un5_async_prescaler_count_cry_9_S, Y => 
        un5_async_prescaler_count_cry_9_Y, FCO => 
        un5_async_prescaler_count_cry_9_Z);
    
    \delay_counter[14]\ : SLE
      port map(D => delay_counter_lm(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(14));
    
    status_dms1_newVal : SLE
      port map(D => drdy_flank_detected_dms1_0_sqmuxa_1_Z, CLK
         => sb_sb_0_FIC_0_CLK, EN => 
        un1_drdy_flank_detected_dms1_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(15));
    
    \spi_tx_data[7]\ : SLE
      port map(D => N_421_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(7));
    
    \delay_counter[0]\ : SLE
      port map(D => delay_counter_lm(0), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(0));
    
    \delay_counter_cry[13]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(13), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(12), S => 
        delay_counter_s(13), Y => delay_counter_cry_Y(13), FCO
         => delay_counter_cry_Z(13));
    
    un1_presetn_inv_i_a3_0_a2_0_x : CFG3
      generic map(INIT => x"10")

      port map(A => sb_sb_0_STAMP_PADDR(3), B => 
        sb_sb_0_STAMP_PADDR(2), C => 
        un1_presetn_inv_i_a3_0_a2_0_1_0_Z, Y => 
        un1_presetn_inv_i_a3_0_a2_0_x_Z);
    
    \dummy[14]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(14), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(14));
    
    \un1_spi_rx_data_0[12]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(12), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(12), Y => N_597);
    
    un1_component_state_9_1 : CFG3
      generic map(INIT => x"FE")

      port map(A => component_state_Z(4), B => 
        component_state_Z(2), C => component_state_Z(0), Y => 
        un1_component_state_9_1_Z);
    
    \delay_counter_cry[7]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(7), C => \GND\, D
         => \GND\, FCI => delay_counter_cry_Z(6), S => 
        delay_counter_s(7), Y => delay_counter_cry_Y(7), FCO => 
        delay_counter_cry_Z(7));
    
    \delay_counter_cry[4]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(4), C => \GND\, D
         => \GND\, FCI => delay_counter_cry_Z(3), S => 
        delay_counter_s(4), Y => delay_counter_cry_Y(4), FCO => 
        delay_counter_cry_Z(4));
    
    \async_prescaler_count[7]\ : SLE
      port map(D => async_prescaler_count_5_Z(7), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(7));
    
    \delay_counter_cry[17]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(17), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(16), S => 
        delay_counter_s(17), Y => delay_counter_cry_Y(17), FCO
         => delay_counter_cry_Z(17));
    
    \async_prescaler_count[6]\ : SLE
      port map(D => async_prescaler_count_5_Z(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(6));
    
    \dummy[26]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(26));
    
    \measurement_dms2[14]\ : SLE
      port map(D => spi_rx_data(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(46));
    
    \delay_counter_lm_0[27]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s_Z(27), Y => 
        delay_counter_lm(27));
    
    un1_request_resync_0_sqmuxa_1_0_0_1 : CFG3
      generic map(INIT => x"7F")

      port map(A => sb_sb_0_STAMP_PADDR(9), B => 
        sb_sb_0_STAMP_PWRITE, C => sb_sb_0_STAMP_PADDR(7), Y => 
        un1_request_resync_0_sqmuxa_1_0_0_1_Z);
    
    \async_prescaler_count[4]\ : SLE
      port map(D => un5_async_prescaler_count_cry_4_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(4));
    
    \delay_counter[13]\ : SLE
      port map(D => delay_counter_lm(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(13));
    
    \delay_counter_RNIKM2J[10]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => delay_counter_Z(11), B => delay_counter_Z(10), 
        C => delay_counter_Z(9), D => delay_counter_Z(8), Y => 
        N_519_i_0_a2_20);
    
    \delay_counter[10]\ : SLE
      port map(D => delay_counter_lm(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(10));
    
    \component_state[5]\ : SLE
      port map(D => component_state_ns(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \GND\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => component_state_Z(5));
    
    un1_request_resync_0_sqmuxa_1_0_0_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => component_state_Z(5), B => config_Z(31), Y
         => N_493);
    
    \un1_spi_rx_data_0[22]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(22), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(22), Y => N_607);
    
    \config[10]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(10), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(10));
    
    \un1_spi_rx_data_0[15]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(15), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(15), Y => N_600);
    
    \PRDATA[17]\ : SLE
      port map(D => N_669, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(17));
    
    \un1_spi_rx_data_2[19]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_638, B => N_604, C => N_107, Y => N_671);
    
    un1_component_state_9_3 : CFG4
      generic map(INIT => x"FFF4")

      port map(A => spi_busy, B => component_state_Z(1), C => 
        spi_enable_1_sqmuxa_1_Z, D => un1_component_state_9_1_Z, 
        Y => un1_component_state_9_3_Z);
    
    \measurement_temp[9]\ : SLE
      port map(D => spi_rx_data(9), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(25));
    
    N_47_i : CFG4
      generic map(INIT => x"F0E0")

      port map(A => sb_sb_0_STAMP_PADDR(5), B => 
        sb_sb_0_STAMP_PADDR(6), C => sb_sb_0_STAMP_PWRITE, D => 
        sb_sb_0_STAMP_PADDR(4), Y => N_47_i_Z);
    
    \spi_request_for[1]\ : SLE
      port map(D => N_570_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_4_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => 
        spi_request_for_Z(1));
    
    \un1_spi_rx_data_2[10]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_629, B => N_595, C => N_107, Y => N_662);
    
    \un1_spi_rx_data_0[17]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(17), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(17), Y => N_602);
    
    \PRDATA[18]\ : SLE
      port map(D => N_670, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(18));
    
    \un1_spi_rx_data_1[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(35), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(3), Y => N_622);
    
    \delay_counter_lm_0[20]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(20), Y => 
        delay_counter_lm(20));
    
    \config[0]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(0));
    
    \dummy[19]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(19));
    
    \un1_spi_rx_data_1[24]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(56), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(24), Y => N_643);
    
    \measurement_dms1[5]\ : SLE
      port map(D => spi_rx_data(5), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(53));
    
    \un1_spi_rx_data_2[31]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_650, B => N_616, C => N_107, Y => N_683);
    
    \measurement_dms2[0]\ : SLE
      port map(D => spi_rx_data(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(32));
    
    \un1_spi_rx_data_0[25]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame\(25), B => config_Z(25), 
        C => sb_sb_0_STAMP_PADDR(8), Y => N_610);
    
    \async_state[0]\ : SLE
      port map(D => N_33_i, CLK => sb_sb_0_FIC_0_CLK, EN => \VCC\, 
        ALn => debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => async_state_Z(0));
    
    un1_drdy_flank_detected_dms1_0_sqmuxa_1_0_0 : CFG3
      generic map(INIT => x"FE")

      port map(A => N_498, B => N_493, C => 
        drdy_flank_detected_dms1_0_sqmuxa_1_Z, Y => 
        un1_drdy_flank_detected_dms1_0_sqmuxa_1_0_0_Z);
    
    \delay_counter_cry[20]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(20), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(19), S => 
        delay_counter_s(20), Y => delay_counter_cry_Y(20), FCO
         => delay_counter_cry_Z(20));
    
    \un1_spi_rx_data_0[27]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame\(27), B => config_Z(27), 
        C => sb_sb_0_STAMP_PADDR(8), Y => N_612);
    
    \measurement_dms2[2]\ : SLE
      port map(D => spi_rx_data(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(34));
    
    \un1_spi_rx_data_1[23]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(55), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(23), Y => N_642);
    
    \un1_spi_rx_data_1[26]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(58), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(26), Y => N_645);
    
    \un1_spi_rx_data[15]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_667, C => 
        spi_rx_data(15), Y => N_700);
    
    \component_state_ns_0_0_0[2]\ : CFG4
      generic map(INIT => x"EFEE")

      port map(A => N_386, B => N_353_i, C => un27_paddr_i_0, D
         => component_state_ns_0_0_0_a3_2_Z(2), Y => 
        component_state_ns(2));
    
    status_dms2_newVal : SLE
      port map(D => drdy_flank_detected_dms2_1_sqmuxa_1, CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_new_avail_0_sqmuxa_3_0_0_Z, 
        ALn => debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(14));
    
    status_temp_overwrittenVal_9 : CFG3
      generic map(INIT => x"04")

      port map(A => N_498, B => \STAMP_0_data_frame\(13), C => 
        N_493, Y => status_temp_overwrittenVal_9_Z);
    
    \un1_spi_rx_data_1[14]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(46), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(14), Y => N_633);
    
    \config[1]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(1));
    
    \un1_spi_rx_data_2_1_1[1]\ : CFG4
      generic map(INIT => x"5553")

      port map(A => \STAMP_0_data_frame\(1), B => 
        \STAMP_0_data_frame\(33), C => sb_sb_0_STAMP_PADDR(9), D
         => sb_sb_0_STAMP_PADDR(7), Y => 
        un1_spi_rx_data_2_1_1_Z(1));
    
    \delay_counter[16]\ : SLE
      port map(D => delay_counter_lm(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(16));
    
    \delay_counter[18]\ : SLE
      port map(D => delay_counter_lm(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(18));
    
    spi_tx_data_0_sqmuxa_RNI8RCF : CFG3
      generic map(INIT => x"C8")

      port map(A => next_state_1_sqmuxa, B => debug_led_net_0, C
         => spi_tx_data_0_sqmuxa_Z, Y => un1_presetn_inv_2_i);
    
    \delay_counter_RNIEFPA[20]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => delay_counter_Z(23), B => delay_counter_Z(22), 
        C => delay_counter_Z(21), D => delay_counter_Z(20), Y => 
        N_519_i_0_a2_14);
    
    \dummy[21]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(21), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(21));
    
    \dummy[16]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(16), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(16));
    
    \component_state_ns_i_a3_i_0_a3_1[4]\ : CFG3
      generic map(INIT => x"80")

      port map(A => next_state_0_sqmuxa_Z, B => N_309, C => 
        component_state_Z(5), Y => N_392);
    
    \async_prescaler_count_5[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => un1_async_prescaler_count, B => 
        un5_async_prescaler_count_cry_6_S, Y => 
        async_prescaler_count_5_Z(6));
    
    spi_dms2_cs_0_sqmuxa : CFG4
      generic map(INIT => x"7F00")

      port map(A => spi_dms2_cs_1_sqmuxa_0_Z, B => N_309, C => 
        config_Z(30), D => component_state_Z(5), Y => 
        spi_dms2_cs_0_sqmuxa_Z);
    
    un5_async_prescaler_count_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(2), C => 
        \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_1_Z, S => 
        un5_async_prescaler_count_cry_2_S, Y => 
        un5_async_prescaler_count_cry_2_Y, FCO => 
        un5_async_prescaler_count_cry_2_Z);
    
    \measurement_dms2[8]\ : SLE
      port map(D => spi_rx_data(8), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(40));
    
    \delay_counter_lm_0[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(26), Y => 
        delay_counter_lm(26));
    
    \un1_spi_rx_data_1[13]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame\(45), B => dummy_Z(13), C
         => sb_sb_0_STAMP_PADDR(8), D => sb_sb_0_STAMP_PADDR(9), 
        Y => N_632);
    
    \un1_spi_rx_data_1[16]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(48), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(16), Y => N_635);
    
    \measurement_dms1[2]\ : SLE
      port map(D => spi_rx_data(2), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(50));
    
    spi_temp_cs_ldmx : CFG4
      generic map(INIT => x"3B31")

      port map(A => spi_temp_cs_0_sqmuxa_Z, B => 
        spi_temp_cs_13_iv, C => config_Z(31), D => 
        \stamp0_spi_temp_cs_c\, Y => spi_temp_cs_ldmx_Z);
    
    \config[23]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(23));
    
    \delay_counter_lm_0[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_332_i, B => N_176, C => delay_counter_s(3), 
        Y => delay_counter_lm(3));
    
    un5_async_prescaler_count_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(3), C => 
        \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_2_Z, S => 
        un5_async_prescaler_count_cry_3_S, Y => 
        un5_async_prescaler_count_cry_3_Y, FCO => 
        un5_async_prescaler_count_cry_3_Z);
    
    \un1_spi_rx_data_2[28]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_647, B => N_613, C => N_107, Y => N_680);
    
    \delay_counter_RNIUVPA[24]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => delay_counter_Z(27), B => delay_counter_Z(26), 
        C => delay_counter_Z(25), D => delay_counter_Z(24), Y => 
        N_519_i_0_a2_16);
    
    \delay_counter[7]\ : SLE
      port map(D => delay_counter_lm(7), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(7));
    
    un1_presetn_inv_i_a3_0_a3_RNIM5LV1 : CFG2
      generic map(INIT => x"E")

      port map(A => un1_presetn_inv_i_a3_0_a3_Z, B => 
        un1_presetn_inv_i_a3_0_a2_0_RNINN9L1_Z, Y => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z);
    
    un1_presetn_inv_i_a3_0_a2_0 : CFG4
      generic map(INIT => x"0001")

      port map(A => sb_sb_0_STAMP_PADDR(6), B => 
        sb_sb_0_STAMP_PADDR(5), C => un1_APBState_1_5, D => 
        un1_presetn_inv_i_a3_0_a2_0_sx_Z, Y => N_486);
    
    \delay_counter_lm_0[15]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(15), Y => 
        delay_counter_lm(15));
    
    \un1_spi_rx_data_1[7]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame\(39), B => dummy_Z(7), C
         => sb_sb_0_STAMP_PADDR(8), D => sb_sb_0_STAMP_PADDR(9), 
        Y => N_626);
    
    \config[19]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(19), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(19));
    
    \config[5]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(5));
    
    \delay_counter_RNIMTFR[4]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => delay_counter_Z(7), B => delay_counter_Z(6), 
        C => delay_counter_Z(5), D => delay_counter_Z(4), Y => 
        N_519_i_0_a2_17);
    
    \component_state_ns_0_0_0_a3_0[2]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => spi_busy, B => component_state_Z(0), C => 
        apb_spi_finished_1_sqmuxa_0, D => N_309, Y => N_386);
    
    next_state_0_sqmuxa : CFG4
      generic map(INIT => x"CCC8")

      port map(A => drdy_flank_detected_dms1_Z, B => config_Z(30), 
        C => drdy_flank_detected_temp_Z, D => 
        drdy_flank_detected_dms2_Z, Y => next_state_0_sqmuxa_Z);
    
    \delay_counter_cry[9]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(9), C => \GND\, D
         => \GND\, FCI => delay_counter_cry_Z(8), S => 
        delay_counter_s(9), Y => delay_counter_cry_Y(9), FCO => 
        delay_counter_cry_Z(9));
    
    spi_temp_cs_0_sqmuxa : CFG4
      generic map(INIT => x"7F00")

      port map(A => un15_delay_counter_Z, B => N_309, C => 
        config_Z(30), D => component_state_Z(5), Y => 
        spi_temp_cs_0_sqmuxa_Z);
    
    measurement_dms1_0_sqmuxa : CFG4
      generic map(INIT => x"0800")

      port map(A => N_309, B => debug_led_net_0, C => spi_busy, D
         => component_state_Z(0), Y => 
        measurement_dms1_0_sqmuxa_Z);
    
    \un1_spi_rx_data_2[21]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_640, B => N_606, C => N_107, Y => N_673);
    
    \PRDATA[24]\ : SLE
      port map(D => N_676, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(24));
    
    un1_presetn_inv_i_a3_0_a2_0_sx : CFG4
      generic map(INIT => x"FFEF")

      port map(A => sb_sb_0_STAMP_PADDR(3), B => 
        sb_sb_0_STAMP_PADDR(2), C => component_state_Z(3), D => 
        sb_sb_0_STAMP_PADDR(4), Y => 
        un1_presetn_inv_i_a3_0_a2_0_sx_Z);
    
    \measurement_temp[13]\ : SLE
      port map(D => spi_rx_data(13), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(29));
    
    \un1_spi_rx_data_2[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_623, B => N_589, C => N_107, Y => N_656);
    
    \spi_tx_data[10]\ : SLE
      port map(D => N_418_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(10));
    
    \status_async_cycles_lm_0[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => status_async_cycles_3_sqmuxa_Z, B => 
        status_async_cycles_s(3), C => 
        status_async_cycles_1_sqmuxa, Y => 
        status_async_cycles_lm(3));
    
    \spi_tx_data_RNO[10]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(10), B => 
        component_state_Z(5), Y => N_418_i);
    
    un1_async_state_0_sqmuxa_0_0_0 : CFG4
      generic map(INIT => x"F2F0")

      port map(A => async_state_Z(0), B => async_state_Z(1), C
         => N_493, D => N_498, Y => un1_async_state_0_sqmuxa_i);
    
    \un1_spi_rx_data_1[30]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(62), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(30), Y => N_649);
    
    drdy_flank_detected_dms2_1_sqmuxa_1_0_a4_0_a3_0 : CFG2
      generic map(INIT => x"8")

      port map(A => component_state_Z(0), B => 
        spi_request_for_Z(0), Y => 
        drdy_flank_detected_dms2_1_sqmuxa_1_0_a4_0_a3_0_Z);
    
    request_resync_1_sqmuxa_1_0_a4 : CFG4
      generic map(INIT => x"0004")

      port map(A => async_state_Z(1), B => async_state_Z(0), C
         => un1_async_prescaler_count, D => 
        un45_async_state_cry_5_Z, Y => request_resync_1_sqmuxa_1);
    
    \measurement_temp[15]\ : SLE
      port map(D => spi_rx_data(15), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(31));
    
    \un1_spi_rx_data[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_655, C => 
        spi_rx_data(3), Y => N_688);
    
    drdy_flank_detected_temp_1_sqmuxa_2_i_0_0 : CFG3
      generic map(INIT => x"FB")

      port map(A => drdy_flank_detected_temp_1_sqmuxa_1, B => 
        stamp0_ready_temp_c, C => N_493, Y => 
        drdy_flank_detected_temp_1_sqmuxa_2_i_0_0_Z);
    
    \dummy[23]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(23), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(23));
    
    \delay_counter_cry[2]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(2), C => \GND\, D
         => \GND\, FCI => delay_counter_cry_Z(1), S => 
        delay_counter_s(2), Y => delay_counter_cry_Y(2), FCO => 
        delay_counter_cry_Z(2));
    
    \async_prescaler_count_5[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => un1_async_prescaler_count, B => 
        un5_async_prescaler_count_s_11_S, Y => 
        async_prescaler_count_5_Z(11));
    
    drdy_flank_detected_dms2_1_sqmuxa_2_i_0_0 : CFG3
      generic map(INIT => x"FB")

      port map(A => drdy_flank_detected_dms2_1_sqmuxa_1, B => 
        stamp0_ready_dms2_c, C => N_493, Y => N_21);
    
    un5_async_prescaler_count_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(5), C => 
        \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_4_Z, S => 
        un5_async_prescaler_count_cry_5_S, Y => 
        un5_async_prescaler_count_cry_5_Y, FCO => 
        un5_async_prescaler_count_cry_5_Z);
    
    \dummy[11]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(11));
    
    \async_prescaler_count_5[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => un1_async_prescaler_count, B => 
        un5_async_prescaler_count_cry_2_S, Y => 
        async_prescaler_count_5_Z(2));
    
    apb_is_atomic_0_sqmuxa_0_a4_i_o3_RNIPU57 : CFG2
      generic map(INIT => x"8")

      port map(A => debug_led_net_0, B => N_353_i, Y => N_178_i);
    
    GND_Z : GND
      port map(Y => \GND\);
    
    \dummy[28]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(28));
    
    \un1_spi_rx_data_2[14]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_633, B => N_599, C => N_107, Y => N_666);
    
    \component_state_ns_0_0_0_a3_2[2]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => apb_spi_finished_Z, B => component_state_Z(3), 
        C => component_state_Z(0), D => N_47_i_Z, Y => 
        component_state_ns_0_0_0_a3_2_Z(2));
    
    \un1_spi_rx_data_2[9]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_628, B => N_107, C => N_594, Y => N_661);
    
    spi_dms1_cs_0_sqmuxa_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => drdy_flank_detected_dms1_Z, B => config_Z(30), 
        C => component_state_Z(5), D => N_309, Y => 
        spi_dms1_cs_0_sqmuxa_3_Z);
    
    \component_state_ns_0_1[0]\ : CFG4
      generic map(INIT => x"F2F0")

      port map(A => component_state_ns_0_a3_0_0_Z(0), B => 
        spi_busy, C => component_state_ns_0_0_Z(0), D => N_309, Y
         => component_state_ns_0_1_Z(0));
    
    un1_component_state_13_0_i_tz : CFG3
      generic map(INIT => x"8C")

      port map(A => un1_component_state_13_0_i_a3_0_1_0_Z, B => 
        N_487, C => component_state_Z(0), Y => N_165_tz);
    
    \async_state_17_iv_0_0_0[1]\ : CFG4
      generic map(INIT => x"FF09")

      port map(A => N_331, B => async_state_Z(1), C => 
        un1_async_state_0_sqmuxa_i, D => 
        request_resync_1_sqmuxa_1, Y => 
        async_state_17_iv_0_0_0_Z(1));
    
    \measurement_temp[0]\ : SLE
      port map(D => spi_rx_data(0), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(16));
    
    \delay_counter_lm_0[11]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(11), Y => 
        delay_counter_lm(11));
    
    \async_state_17_iv_0_0_a2[1]\ : CFG4
      generic map(INIT => x"0010")

      port map(A => spi_request_for_Z(1), B => async_state_Z(1), 
        C => N_309, D => spi_busy, Y => N_499);
    
    \measurement_temp[1]\ : SLE
      port map(D => spi_rx_data(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(17));
    
    \dummy[5]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(5), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(5));
    
    \component_state_ns_i_a3_i_0[4]\ : CFG4
      generic map(INIT => x"FFF2")

      port map(A => component_state_Z(1), B => spi_busy, C => 
        N_392, D => next_state_1_sqmuxa, Y => N_28);
    
    \spi_tx_data[0]\ : SLE
      port map(D => N_428_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(0));
    
    \spi_tx_data[14]\ : SLE
      port map(D => N_414_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(14));
    
    \un1_spi_rx_data_0[31]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame\(31), B => config_Z(31), 
        C => sb_sb_0_STAMP_PADDR(8), Y => N_616);
    
    un5_async_prescaler_count_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(6), C => 
        \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_5_Z, S => 
        un5_async_prescaler_count_cry_6_S, Y => 
        un5_async_prescaler_count_cry_6_Y, FCO => 
        un5_async_prescaler_count_cry_6_Z);
    
    \measurement_temp[12]\ : SLE
      port map(D => spi_rx_data(12), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(28));
    
    \un1_spi_rx_data_2[13]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_632, B => N_107, C => N_598, Y => N_665);
    
    \un1_spi_rx_data[7]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_659, C => 
        spi_rx_data(7), Y => un1_spi_rx_data_Z(7));
    
    \PRDATA[20]\ : SLE
      port map(D => N_672, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(20));
    
    \delay_counter_cry[3]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(3), C => \GND\, D
         => \GND\, FCI => delay_counter_cry_Z(2), S => 
        delay_counter_s(3), Y => delay_counter_cry_Y(3), FCO => 
        delay_counter_cry_Z(3));
    
    \async_state_RNO[0]\ : CFG4
      generic map(INIT => x"0012")

      port map(A => N_275, B => un1_async_state_0_sqmuxa_i, C => 
        async_state_Z(0), D => request_resync_1_sqmuxa_1, Y => 
        N_33_i);
    
    \un1_spi_rx_data_2[16]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_635, B => N_601, C => N_107, Y => N_668);
    
    \delay_counter_RNIG01L3[10]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_519_i_0_a2_14, B => N_519_i_0_a2_25, C => 
        N_519_i_0_a2_20, D => N_519_i_0_a2_15, Y => N_309);
    
    \un1_spi_rx_data[6]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_658, C => 
        spi_rx_data(6), Y => un1_spi_rx_data_Z(6));
    
    \un1_spi_rx_data_2[1]\ : CFG4
      generic map(INIT => x"B133")

      port map(A => sb_sb_0_STAMP_PADDR(8), B => 
        un1_spi_rx_data_2_1_1_Z(1), C => dummy_Z(1), D => 
        sb_sb_0_STAMP_PADDR(9), Y => N_653);
    
    drdy_flank_detected_dms2_RNO : CFG1
      generic map(INIT => "01")

      port map(A => stamp0_ready_dms2_c, Y => 
        stamp0_ready_dms2_c_i);
    
    un5_async_prescaler_count_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(8), C => 
        \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_cry_7_Z, S => 
        un5_async_prescaler_count_cry_8_S, Y => 
        un5_async_prescaler_count_cry_8_Y, FCO => 
        un5_async_prescaler_count_cry_8_Z);
    
    \dummy[9]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(9));
    
    \delay_counter_cry[25]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(25), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(24), S => 
        delay_counter_s(25), Y => delay_counter_cry_Y(25), FCO
         => delay_counter_cry_Z(25));
    
    un1_component_state_14_0_i_o2_RNO : CFG4
      generic map(INIT => x"70F0")

      port map(A => drdy_flank_detected_dms1_Z, B => config_Z(30), 
        C => component_state_Z(5), D => N_309, Y => spi_N_5_mux_i);
    
    \PRDATA[23]\ : SLE
      port map(D => N_675, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(23));
    
    apb_is_atomic_0_sqmuxa_0_a4_i_o3 : CFG2
      generic map(INIT => x"8")

      port map(A => sb_sb_0_STAMP_PENABLE, B => 
        component_state_Z(4), Y => N_353_i);
    
    \delay_counter_cry[8]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(8), C => \GND\, D
         => \GND\, FCI => delay_counter_cry_Z(7), S => 
        delay_counter_s(8), Y => delay_counter_cry_Y(8), FCO => 
        delay_counter_cry_Z(8));
    
    \un1_spi_rx_data[5]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_657, C => 
        spi_rx_data(5), Y => N_690);
    
    \measurement_dms1[3]\ : SLE
      port map(D => spi_rx_data(3), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(51));
    
    un1_presetn_inv_i_a3_0_a2_0_RNINN9L1 : CFG4
      generic map(INIT => x"8000")

      port map(A => N_486, B => PRDATA_684_1_Z, C => 
        debug_led_net_0, D => un1_spi_rx_data_sn_N_5, Y => 
        un1_presetn_inv_i_a3_0_a2_0_RNINN9L1_Z);
    
    status_temp_overwrittenVal : SLE
      port map(D => status_temp_overwrittenVal_9_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_new_avail_0_sqmuxa_2_0_0_Z, 
        ALn => debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, 
        SD => \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(10));
    
    \delay_counter_lm_0[0]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => delay_counter_cry_Y(0), B => 
        apb_spi_finished_0_sqmuxa_1, C => N_176, Y => 
        delay_counter_lm(0));
    
    \delay_counter_cry[26]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(26), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(25), S => 
        delay_counter_s(26), Y => delay_counter_cry_Y(26), FCO
         => delay_counter_cry_Z(26));
    
    \async_prescaler_count[8]\ : SLE
      port map(D => async_prescaler_count_5_Z(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(8));
    
    \measurement_dms1[1]\ : SLE
      port map(D => spi_rx_data(1), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(49));
    
    \async_state_RNO_0[0]\ : CFG4
      generic map(INIT => x"0301")

      port map(A => component_state_Z(0), B => 
        component_state_Z(5), C => N_318, D => N_499, Y => N_275);
    
    \spi_tx_data[12]\ : SLE
      port map(D => N_416_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(12));
    
    \delay_counter[27]\ : SLE
      port map(D => delay_counter_lm(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(27));
    
    \un1_spi_rx_data_0[19]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(19), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(19), Y => N_604);
    
    drdy_flank_detected_dms2_1_sqmuxa_1_0_a4_0_a3 : CFG4
      generic map(INIT => x"1000")

      port map(A => spi_request_for_Z(1), B => spi_busy, C => 
        drdy_flank_detected_dms2_1_sqmuxa_1_0_a4_0_a3_0_Z, D => 
        N_309, Y => drdy_flank_detected_dms2_1_sqmuxa_1);
    
    \config[22]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(22));
    
    \PRDATA[30]\ : SLE
      port map(D => N_682, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(30));
    
    \un1_spi_rx_data_0[10]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(10), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(10), Y => N_595);
    
    \PRDATA[11]\ : SLE
      port map(D => un1_spi_rx_data_Z(11), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_presetn_inv_i_a3_0_a3_Z, ALn
         => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => sb_sb_0_STAMP_PRDATA(11));
    
    \spi_tx_data_RNO[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(5), B => 
        component_state_Z(5), Y => N_423_i);
    
    \un1_spi_rx_data[11]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_663, C => 
        spi_rx_data(11), Y => un1_spi_rx_data_Z(11));
    
    status_dms1_overwrittenVal : SLE
      port map(D => N_270_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_drdy_flank_detected_dms1_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(12));
    
    \measurement_temp[14]\ : SLE
      port map(D => spi_rx_data(14), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_temp_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(30));
    
    \dummy[13]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(13), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(13));
    
    \config[8]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(8));
    
    \measurement_dms1[10]\ : SLE
      port map(D => spi_rx_data(10), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(58));
    
    \component_state_RNIE2K05[3]\ : CFG4
      generic map(INIT => x"2A0A")

      port map(A => delay_counterlde_0_0_a3_2, B => N_309, C => 
        component_state_Z(3), D => component_state_Z(5), Y => 
        N_381);
    
    \config[6]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(6), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(6));
    
    \status_async_cycles_lm_0[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => status_async_cycles_3_sqmuxa_Z, B => 
        status_async_cycles_s(4), C => 
        status_async_cycles_1_sqmuxa, Y => 
        status_async_cycles_lm(4));
    
    spi_request_for_2_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => un15_delay_counter_Z, B => N_309, C => 
        config_Z(30), D => component_state_Z(5), Y => 
        spi_request_for_2_sqmuxa_Z);
    
    un1_component_state_17_0_i_a3_0 : CFG4
      generic map(INIT => x"0040")

      port map(A => spi_request_for_Z(1), B => 
        spi_request_for_Z(0), C => N_309, D => spi_busy, Y => 
        un1_component_state_17_0_i_a3_0_Z);
    
    \dummy[8]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(8));
    
    spi_dms2_cs_13_iv_i : CFG3
      generic map(INIT => x"13")

      port map(A => component_state_Z(3), B => 
        spi_dms2_cs_1_sqmuxa_1_Z, C => sb_sb_0_STAMP_PADDR(5), Y
         => spi_dms2_cs_13_iv_i_Z);
    
    \measurement_dms1[4]\ : SLE
      port map(D => spi_rx_data(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(52));
    
    \measurement_dms1[11]\ : SLE
      port map(D => spi_rx_data(11), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(59));
    
    \un1_spi_rx_data[13]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_665, C => 
        spi_rx_data(13), Y => N_698);
    
    \un1_spi_rx_data_1[9]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame\(41), B => dummy_Z(9), C
         => sb_sb_0_STAMP_PADDR(8), D => sb_sb_0_STAMP_PADDR(9), 
        Y => N_628);
    
    \component_state_RNO[0]\ : CFG4
      generic map(INIT => x"AF88")

      port map(A => spi_busy, B => component_state_Z(1), C => 
        N_309, D => component_state_Z(0), Y => N_151_i);
    
    \delay_counter_cry[18]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(18), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(17), S => 
        delay_counter_s(18), Y => delay_counter_cry_Y(18), FCO
         => delay_counter_cry_Z(18));
    
    \delay_counter_cry[24]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(24), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(23), S => 
        delay_counter_s(24), Y => delay_counter_cry_Y(24), FCO
         => delay_counter_cry_Z(24));
    
    \dummy[18]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(18), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(18));
    
    \un1_spi_rx_data_0[29]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \STAMP_0_data_frame\(29), B => config_Z(29), 
        C => sb_sb_0_STAMP_PADDR(8), Y => N_614);
    
    \status_async_cycles[2]\ : SLE
      port map(D => status_async_cycles_lm(2), CLK => 
        sb_sb_0_FIC_0_CLK, EN => status_async_cyclese, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(5));
    
    un1_spi_rx_data_sn_m4 : CFG2
      generic map(INIT => x"1")

      port map(A => sb_sb_0_STAMP_PADDR(8), B => 
        sb_sb_0_STAMP_PADDR(9), Y => un1_spi_rx_data_sn_N_5);
    
    \delay_counter_cry[22]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(22), C => \GND\, 
        D => \GND\, FCI => delay_counter_cry_Z(21), S => 
        delay_counter_s(22), Y => delay_counter_cry_Y(22), FCO
         => delay_counter_cry_Z(22));
    
    \un1_spi_rx_data_1[8]\ : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \STAMP_0_data_frame\(40), B => dummy_Z(8), C
         => sb_sb_0_STAMP_PADDR(8), D => sb_sb_0_STAMP_PADDR(9), 
        Y => N_627);
    
    \un1_spi_rx_data_0[20]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(20), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(20), Y => N_605);
    
    \spi_request_for_RNO[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => spi_dms2_cs_1_sqmuxa_1_Z, B => 
        component_state_Z(3), Y => N_569_i);
    
    \async_state_17_iv_0_0[1]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => async_state_17_iv_0_0_a3_0_1_Z(1), B => N_499, 
        C => un1_async_state_0_sqmuxa_i, D => 
        async_state_17_iv_0_0_0_Z(1), Y => async_state_17(1));
    
    spi_tx_data_0_sqmuxa : CFG3
      generic map(INIT => x"80")

      port map(A => config_Z(30), B => component_state_Z(5), C
         => N_309, Y => spi_tx_data_0_sqmuxa_Z);
    
    \async_prescaler_count[5]\ : SLE
      port map(D => un5_async_prescaler_count_cry_5_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(5));
    
    \un1_spi_rx_data_2[22]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_641, B => N_607, C => N_107, Y => N_674);
    
    spi_temp_cs_13_iv_0_0_0 : CFG3
      generic map(INIT => x"EC")

      port map(A => component_state_Z(3), B => 
        spi_request_for_2_sqmuxa_Z, C => sb_sb_0_STAMP_PADDR(6), 
        Y => spi_temp_cs_13_iv);
    
    \spi_tx_data[4]\ : SLE
      port map(D => N_424_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(4));
    
    \delay_counter_cry[5]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => \VCC\, B => delay_counter_Z(5), C => \GND\, D
         => \GND\, FCI => delay_counter_cry_Z(4), S => 
        delay_counter_s(5), Y => delay_counter_cry_Y(5), FCO => 
        delay_counter_cry_Z(5));
    
    \config[26]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(26), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(26));
    
    \un1_spi_rx_data_1[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(36), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(4), Y => N_623);
    
    \PRDATA[25]\ : SLE
      port map(D => N_677, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(25));
    
    \spi_tx_data_RNO[4]\ : CFG2
      generic map(INIT => x"E")

      port map(A => sb_sb_0_STAMP_PWDATA(4), B => 
        component_state_Z(5), Y => N_424_i);
    
    \delay_counter_lm_0[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(2), Y => 
        delay_counter_lm(2));
    
    \status_async_cycles[0]\ : SLE
      port map(D => status_async_cycles_lm(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => status_async_cyclese, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(3));
    
    un45_async_state_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => config_Z(27), B => \STAMP_0_data_frame\(6), C
         => \GND\, D => \GND\, FCI => un45_async_state_cry_2_Z, S
         => un45_async_state_cry_3_S, Y => 
        un45_async_state_cry_3_Y, FCO => un45_async_state_cry_3_Z);
    
    request_resync_1_sqmuxa_2_i_0_0 : CFG2
      generic map(INIT => x"E")

      port map(A => request_resync_1_sqmuxa_1, B => N_493, Y => 
        N_40);
    
    \delay_counter_lm_0[23]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(23), Y => 
        delay_counter_lm(23));
    
    \PRDATA[0]\ : SLE
      port map(D => N_685, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_Z, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_STAMP_PRDATA(0));
    
    \delay_counter_RNI20MA[16]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => delay_counter_Z(19), B => delay_counter_Z(18), 
        C => delay_counter_Z(17), D => delay_counter_Z(16), Y => 
        N_519_i_0_a2_15);
    
    un1_component_state_14_0_i_o2 : CFG2
      generic map(INIT => x"D")

      port map(A => spi_N_5_mux_i, B => config_Z(31), Y => N_279);
    
    \un1_spi_rx_data_2[25]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_644, B => N_610, C => N_107, Y => N_677);
    
    un1_presetn_inv_i_a3_0_a3 : CFG4
      generic map(INIT => x"0800")

      port map(A => N_486, B => debug_led_net_0, C => 
        sb_sb_0_STAMP_PWRITE, D => N_319, Y => 
        un1_presetn_inv_i_a3_0_a3_Z);
    
    un1_component_state_14_0_i : CFG4
      generic map(INIT => x"D000")

      port map(A => component_state_Z(0), B => 
        un1_component_state_14_0_i_a3_0_s_0_Z, C => N_279, D => 
        N_487, Y => N_167);
    
    \status_async_cycles[3]\ : SLE
      port map(D => status_async_cycles_lm(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => status_async_cyclese, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => \STAMP_0_data_frame\(6));
    
    \delay_counter_lm_0[12]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(12), Y => 
        delay_counter_lm(12));
    
    \async_prescaler_count[3]\ : SLE
      port map(D => un5_async_prescaler_count_cry_3_S, CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(3));
    
    \spi_tx_data[5]\ : SLE
      port map(D => N_423_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(5));
    
    \un1_spi_rx_data_2[27]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_646, B => N_612, C => N_107, Y => N_679);
    
    \measurement_dms1[6]\ : SLE
      port map(D => spi_rx_data(6), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms1_0_sqmuxa_1_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(54));
    
    un1_presetn_inv_i_a3_0_a2_0_RNINN9L1_0 : CFG1
      generic map(INIT => "01")

      port map(A => un1_presetn_inv_i_a3_0_a2_0_RNINN9L1_Z, Y => 
        N_1454_i);
    
    status_async_cycles_s_831 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => \STAMP_0_data_frame\(3), C => 
        \GND\, D => \GND\, FCI => \VCC\, S => 
        status_async_cycles_s_831_S, Y => 
        status_async_cycles_s_831_Y, FCO => 
        status_async_cycles_s_831_FCO);
    
    \un1_spi_rx_data[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_652, B => un1_spi_rx_data_sn_N_5, C => 
        spi_rx_data(0), Y => N_685);
    
    \delay_counter_RNICQEC2[12]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_519_i_0_a2_19, B => N_519_i_0_a2_18, C => 
        N_519_i_0_a2_17, D => N_519_i_0_a2_16, Y => 
        N_519_i_0_a2_25);
    
    \dummy[22]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(22), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(22));
    
    apb_spi_finished_1_sqmuxa_0_0 : CFG2
      generic map(INIT => x"8")

      port map(A => spi_request_for_Z(1), B => 
        spi_request_for_Z(0), Y => apb_spi_finished_1_sqmuxa_0);
    
    drdy_flank_detected_dms1 : SLE
      port map(D => stamp0_ready_dms1_c_i, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_23, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => drdy_flank_detected_dms1_Z);
    
    \PRDATA[9]\ : SLE
      port map(D => un1_spi_rx_data_Z(9), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_presetn_inv_i_a3_0_a3_Z, ALn
         => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => sb_sb_0_STAMP_PRDATA(9));
    
    un1_spi_rx_data_sn_m3_0_m2 : CFG3
      generic map(INIT => x"A3")

      port map(A => sb_sb_0_STAMP_PADDR(8), B => 
        sb_sb_0_STAMP_PADDR(7), C => sb_sb_0_STAMP_PADDR(9), Y
         => N_107);
    
    \delay_counter_lm_0[9]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(9), Y => 
        delay_counter_lm(9));
    
    \PRDATA[8]\ : SLE
      port map(D => un1_spi_rx_data_Z(8), CLK => 
        sb_sb_0_FIC_0_CLK, EN => un1_presetn_inv_i_a3_0_a3_Z, ALn
         => \VCC\, ADn => \VCC\, SLn => \VCC\, SD => \GND\, LAT
         => \GND\, Q => sb_sb_0_STAMP_PRDATA(8));
    
    \un1_spi_rx_data_1[28]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(60), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(28), Y => N_647);
    
    \delay_counter[4]\ : SLE
      port map(D => delay_counter_lm(4), CLK => sb_sb_0_FIC_0_CLK, 
        EN => delay_countere, ALn => debug_led_net_0_arst, ADn
         => \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        delay_counter_Z(4));
    
    status_async_cycles_1_sqmuxa_0_a2_0_a3 : CFG3
      generic map(INIT => x"02")

      port map(A => async_state_Z(0), B => async_state_Z(1), C
         => un1_async_prescaler_count, Y => 
        status_async_cycles_1_sqmuxa);
    
    \dummy[3]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(3), CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        un1_request_resync_0_sqmuxa_1_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => N_103_i, SD
         => \GND\, LAT => \GND\, Q => dummy_Z(3));
    
    \spi_tx_data[9]\ : SLE
      port map(D => N_419_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(9));
    
    un1_presetn_inv_i_a3_0_a2_0_1_0 : CFG4
      generic map(INIT => x"0002")

      port map(A => component_state_Z(3), B => 
        sb_sb_0_STAMP_PADDR(4), C => sb_sb_0_STAMP_PADDR(5), D
         => sb_sb_0_STAMP_PADDR(6), Y => 
        un1_presetn_inv_i_a3_0_a2_0_1_0_Z);
    
    \un1_spi_rx_data[9]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_661, C => 
        spi_rx_data(9), Y => un1_spi_rx_data_Z(9));
    
    \PRDATA[22]\ : SLE
      port map(D => N_674, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(22));
    
    \status_async_cycles_lm_0[5]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => status_async_cycles_3_sqmuxa_Z, B => 
        status_async_cycles_s_Z(5), C => 
        status_async_cycles_1_sqmuxa, Y => 
        status_async_cycles_lm(5));
    
    \un1_spi_rx_data_2_1_1[2]\ : CFG4
      generic map(INIT => x"5553")

      port map(A => \STAMP_0_data_frame\(2), B => 
        \STAMP_0_data_frame\(34), C => sb_sb_0_STAMP_PADDR(9), D
         => sb_sb_0_STAMP_PADDR(7), Y => 
        un1_spi_rx_data_2_1_1_Z(2));
    
    \PRDATA[29]\ : SLE
      port map(D => N_681, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_RNIM5LV1_Z, ALn => \VCC\, ADn
         => \VCC\, SLn => N_1454_i, SD => \GND\, LAT => \GND\, Q
         => sb_sb_0_STAMP_PRDATA(29));
    
    \status_async_cycles_lm_0[0]\ : CFG4
      generic map(INIT => x"33FA")

      port map(A => status_async_cycles_2_sqmuxa_Z, B => 
        \STAMP_0_data_frame\(3), C => 
        status_async_cycles_3_sqmuxa_Z, D => 
        status_async_cycles_1_sqmuxa, Y => 
        status_async_cycles_lm(0));
    
    \delay_counter_lm_0[14]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(14), Y => 
        delay_counter_lm(14));
    
    \async_prescaler_count[0]\ : SLE
      port map(D => async_prescaler_count_5_Z(0), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => async_prescaler_count_Z(0));
    
    spi_dms2_cs : SLE
      port map(D => spi_dms2_cs_13_iv_i_Z, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_162, ALn => 
        debug_led_net_0_arst, ADn => \GND\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => stamp0_spi_dms2_cs_c);
    
    \delay_counter[17]\ : SLE
      port map(D => delay_counter_lm(17), CLK => 
        sb_sb_0_FIC_0_CLK, EN => delay_countere, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => delay_counter_Z(17));
    
    \async_prescaler_count_5[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => un1_async_prescaler_count, B => 
        un5_async_prescaler_count_cry_8_S, Y => 
        async_prescaler_count_5_Z(8));
    
    \un1_spi_rx_data_2[0]\ : CFG4
      generic map(INIT => x"B133")

      port map(A => sb_sb_0_STAMP_PADDR(8), B => 
        un1_spi_rx_data_2_1_1_Z(0), C => dummy_Z(0), D => 
        sb_sb_0_STAMP_PADDR(9), Y => N_652);
    
    \status_async_cycles_s[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => \STAMP_0_data_frame\(8), C => 
        \GND\, D => \GND\, FCI => status_async_cycles_cry_Z(4), S
         => status_async_cycles_s_Z(5), Y => 
        status_async_cycles_s_Y(5), FCO => 
        status_async_cycles_s_FCO(5));
    
    \component_state_ns_0_a3_0_0[0]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => spi_request_for_Z(1), B => 
        component_state_Z(0), C => spi_request_for_Z(0), Y => 
        component_state_ns_0_a3_0_0_Z(0));
    
    \config_RNO[31]\ : CFG2
      generic map(INIT => x"2")

      port map(A => sb_sb_0_STAMP_PWDATA(31), B => 
        component_state_Z(5), Y => N_266_i);
    
    \un1_spi_rx_data_1[21]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(53), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(21), Y => N_640);
    
    \config[27]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(27), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(27));
    
    PRDATA_684_1 : CFG4
      generic map(INIT => x"0D06")

      port map(A => sb_sb_0_STAMP_PADDR(9), B => 
        sb_sb_0_STAMP_PADDR(8), C => sb_sb_0_STAMP_PWRITE, D => 
        sb_sb_0_STAMP_PADDR(7), Y => PRDATA_684_1_Z);
    
    \config[28]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(28), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(28));
    
    \component_state[4]\ : SLE
      port map(D => component_state_ns(1), CLK => 
        sb_sb_0_FIC_0_CLK, EN => \VCC\, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => component_state_Z(4));
    
    \un1_spi_rx_data_1[18]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(50), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(18), Y => N_637);
    
    \component_state_RNIT8HJ[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => spi_busy, B => component_state_Z(1), Y => 
        N_332_i);
    
    spi_enable_RNO_0 : CFG4
      generic map(INIT => x"0703")

      port map(A => apb_spi_finished_Z, B => component_state_Z(3), 
        C => un1_component_state_9_3_Z, D => N_47_i_Z, Y => 
        un1_component_state_9_i);
    
    drdy_flank_detected_dms1_0_sqmuxa_1 : CFG4
      generic map(INIT => x"0800")

      port map(A => un3_spi_busy, B => N_309, C => spi_busy, D
         => component_state_Z(0), Y => 
        drdy_flank_detected_dms1_0_sqmuxa_1_Z);
    
    \async_state_17_iv_0_0_o2_RNIPJEP5[1]\ : CFG3
      generic map(INIT => x"AB")

      port map(A => N_381, B => spi_busy, C => N_318, Y => 
        delay_counterlde_0_0_0);
    
    \un1_spi_rx_data_0[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \STAMP_0_data_frame\(3), B => 
        sb_sb_0_STAMP_PADDR(8), C => config_Z(3), Y => N_588);
    
    \component_state[0]\ : SLE
      port map(D => N_151_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        \VCC\, ALn => debug_led_net_0_arst, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => 
        component_state_Z(0));
    
    \measurement_dms2[4]\ : SLE
      port map(D => spi_rx_data(4), CLK => sb_sb_0_FIC_0_CLK, EN
         => measurement_dms2_1_sqmuxa_Z, ALn => \VCC\, ADn => 
        \VCC\, SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        \STAMP_0_data_frame\(36));
    
    un5_async_prescaler_count_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => \VCC\, B => async_prescaler_count_Z(1), C => 
        \GND\, D => \GND\, FCI => 
        un5_async_prescaler_count_s_1_837_FCO, S => 
        un5_async_prescaler_count_cry_1_S, Y => 
        un5_async_prescaler_count_cry_1_Y, FCO => 
        un5_async_prescaler_count_cry_1_Z);
    
    \config[24]\ : SLE
      port map(D => sb_sb_0_STAMP_PWDATA(24), CLK => 
        sb_sb_0_FIC_0_CLK, EN => config_143, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => config_Z(24));
    
    \spi_tx_data[8]\ : SLE
      port map(D => N_420_i, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_2_i, ALn => \VCC\, ADn => \VCC\, SLn => 
        \VCC\, SD => \GND\, LAT => \GND\, Q => spi_tx_data_Z(8));
    
    drdy_flank_detected_temp : SLE
      port map(D => stamp0_ready_temp_c_i, CLK => 
        sb_sb_0_FIC_0_CLK, EN => 
        drdy_flank_detected_temp_1_sqmuxa_2_i_0_0_Z, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => drdy_flank_detected_temp_Z);
    
    \un1_spi_rx_data[10]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un1_spi_rx_data_sn_N_5, B => N_662, C => 
        spi_rx_data(10), Y => un1_spi_rx_data_Z(10));
    
    \un1_spi_rx_data_2[2]\ : CFG4
      generic map(INIT => x"B133")

      port map(A => sb_sb_0_STAMP_PADDR(8), B => 
        un1_spi_rx_data_2_1_1_Z(2), C => dummy_Z(2), D => 
        sb_sb_0_STAMP_PADDR(9), Y => N_654);
    
    \PRDATA[4]\ : SLE
      port map(D => N_689, CLK => sb_sb_0_FIC_0_CLK, EN => 
        un1_presetn_inv_i_a3_0_a3_Z, ALn => \VCC\, ADn => \VCC\, 
        SLn => \VCC\, SD => \GND\, LAT => \GND\, Q => 
        sb_sb_0_STAMP_PRDATA(4));
    
    drdy_flank_detected_dms2 : SLE
      port map(D => stamp0_ready_dms2_c_i, CLK => 
        sb_sb_0_FIC_0_CLK, EN => N_21, ALn => 
        debug_led_net_0_arst, ADn => \VCC\, SLn => \VCC\, SD => 
        \GND\, LAT => \GND\, Q => drdy_flank_detected_dms2_Z);
    
    \delay_counter_lm_0[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_176, B => delay_counter_s(5), Y => 
        delay_counter_lm(5));
    
    \un1_spi_rx_data_1[11]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \STAMP_0_data_frame\(43), B => 
        sb_sb_0_STAMP_PADDR(9), C => dummy_Z(11), Y => N_630);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity sb is

    port( DAPI_RX            : in    std_logic;
          DEVRST_N           : in    std_logic;
          MISO               : in    std_logic;
          RXSM_LO            : in    std_logic;
          RXSM_SODS          : in    std_logic;
          RXSM_SOE           : in    std_logic;
          TM_RX              : in    std_logic;
          stamp0_ready_dms1  : in    std_logic;
          stamp0_ready_dms2  : in    std_logic;
          stamp0_ready_temp  : in    std_logic;
          stamp0_spi_miso    : in    std_logic;
          DAPI_TX            : out   std_logic;
          GPIO_6_M2F         : out   std_logic;
          LED_HEARTBEAT      : out   std_logic;
          LED_RECORDING      : out   std_logic;
          MOSI               : out   std_logic;
          SCLK               : out   std_logic;
          TM_TX              : out   std_logic;
          adc_clk            : out   std_logic;
          adc_start          : out   std_logic;
          debug_led          : out   std_logic;
          nCS1               : out   std_logic;
          nCS2               : out   std_logic;
          resetn             : out   std_logic;
          stamp0_spi_clock   : out   std_logic;
          stamp0_spi_dms1_cs : out   std_logic;
          stamp0_spi_dms2_cs : out   std_logic;
          stamp0_spi_mosi    : out   std_logic;
          stamp0_spi_temp_cs : out   std_logic
        );

end sb;

architecture DEF_ARCH of sb is 

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component TRIBUFF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component Memory
    port( sb_sb_0_STAMP_PADDR   : in    std_logic_vector(11 downto 0) := (others => 'U');
          dataReady_0           : in    std_logic := 'U';
          STAMP_0_data_frame    : in    std_logic_vector(63 downto 0) := (others => 'U');
          sb_sb_0_Memory_PRDATA : out   std_logic_vector(31 downto 0);
          sb_sb_0_STAMP_PWDATA  : in    std_logic_vector(31 downto 0) := (others => 'U');
          nCS1_c                : out   std_logic;
          nCS2_c                : out   std_logic;
          MISO_c                : in    std_logic := 'U';
          SCLK_c                : out   std_logic;
          mosi_1                : out   std_logic;
          mosi_cl               : out   std_logic;
          sb_sb_0_STAMP_PENABLE : in    std_logic := 'U';
          sb_sb_0_STAMP_PWRITE  : in    std_logic := 'U';
          sb_sb_0_Memory_PSELx  : in    std_logic := 'U';
          un1_APBState_1_5_1z   : out   std_logic;
          resetn                : in    std_logic := 'U';
          sb_sb_0_Memory_PREADY : out   std_logic;
          GPIO_6_M2F_c          : in    std_logic := 'U';
          sb_sb_0_FIC_0_CLK     : in    std_logic := 'U';
          resetn_arst           : in    std_logic := 'U'
        );
  end component;

  component sb_sb
    port( sb_sb_0_STAMP_PADDR      : out   std_logic_vector(11 downto 0);
          sb_sb_0_STAMP_PWDATA     : out   std_logic_vector(31 downto 0);
          dataReady_0              : in    std_logic := 'U';
          sb_sb_0_Memory_PRDATA    : in    std_logic_vector(31 downto 0) := (others => 'U');
          sb_sb_0_STAMP_PRDATA     : in    std_logic_vector(31 downto 0) := (others => 'U');
          TM_TX                    : out   std_logic;
          TM_RX                    : in    std_logic := 'U';
          DAPI_TX                  : out   std_logic;
          DAPI_RX                  : in    std_logic := 'U';
          sb_sb_0_GPIO_3_M2F       : out   std_logic;
          sb_sb_0_GPIO_4_M2F       : out   std_logic;
          sb_sb_0_STAMP_PENABLE    : out   std_logic;
          sb_sb_0_STAMP_PWRITE     : out   std_logic;
          LED_HEARTBEAT_c          : out   std_logic;
          LED_RECORDING_c          : out   std_logic;
          GPIO_6_M2F_c             : out   std_logic;
          RXSM_LO_c                : in    std_logic := 'U';
          RXSM_SOE_c               : in    std_logic := 'U';
          RXSM_SODS_c              : in    std_logic := 'U';
          sb_sb_0_Memory_PSELx     : out   std_logic;
          sb_sb_0_STAMP_PSELx      : out   std_logic;
          sb_sb_0_Memory_PREADY    : in    std_logic := 'U';
          sb_sb_0_STAMP_PREADY     : in    std_logic := 'U';
          sb_sb_0_FIC_0_CLK        : out   std_logic;
          adc_clk_c                : out   std_logic;
          DEVRST_N                 : in    std_logic := 'U';
          sb_sb_0_POWER_ON_RESET_N : out   std_logic
        );
  end component;

  component STAMP
    port( sb_sb_0_STAMP_PADDR   : in    std_logic_vector(11 downto 2) := (others => 'U');
          STAMP_0_data_frame    : out   std_logic_vector(63 downto 0);
          sb_sb_0_STAMP_PRDATA  : out   std_logic_vector(31 downto 0);
          dataReady_0           : out   std_logic;
          sb_sb_0_STAMP_PWDATA  : in    std_logic_vector(31 downto 0) := (others => 'U');
          stamp0_spi_miso_c     : in    std_logic := 'U';
          stamp0_spi_clock_c    : out   std_logic;
          mosi_1_0              : out   std_logic;
          mosi_cl_0             : out   std_logic;
          sb_sb_0_STAMP_PSELx   : in    std_logic := 'U';
          sb_sb_0_STAMP_PENABLE : in    std_logic := 'U';
          un1_APBState_1_5      : in    std_logic := 'U';
          sb_sb_0_STAMP_PWRITE  : in    std_logic := 'U';
          sb_sb_0_STAMP_PREADY  : out   std_logic;
          debug_led_net_0       : in    std_logic := 'U';
          stamp0_spi_dms1_cs_c  : out   std_logic;
          stamp0_spi_temp_cs_c  : out   std_logic;
          stamp0_spi_dms2_cs_c  : out   std_logic;
          sb_sb_0_FIC_0_CLK     : in    std_logic := 'U';
          debug_led_net_0_arst  : in    std_logic := 'U';
          stamp0_ready_dms1_c   : in    std_logic := 'U';
          stamp0_ready_temp_c   : in    std_logic := 'U';
          stamp0_ready_dms2_c   : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal STAMP_0_data_frame : std_logic_vector(63 downto 0);
    signal \Memory_0.dataReady\ : std_logic_vector(0 to 0);
    signal sb_sb_0_STAMP_PADDR : std_logic_vector(11 downto 0);
    signal sb_sb_0_Memory_PRDATA : std_logic_vector(31 downto 0);
    signal sb_sb_0_STAMP_PRDATA : std_logic_vector(31 downto 0);
    signal sb_sb_0_STAMP_PWDATA : std_logic_vector(31 downto 0);
    signal \GND\, sb_sb_0_GPIO_3_M2F, sb_sb_0_FIC_0_CLK, 
        sb_sb_0_STAMP_PENABLE, sb_sb_0_STAMP_PWRITE, 
        sb_sb_0_Memory_PREADY, sb_sb_0_POWER_ON_RESET_N, 
        sb_sb_0_GPIO_4_M2F, \VCC\, sb_sb_0_STAMP_PREADY, 
        sb_sb_0_STAMP_PSELx, mosi_1, mosi_1_0, 
        debug_led_net_0_arst, resetn_arst, NN_1, debug_led_net_0, 
        sb_sb_0_Memory_PSELx, MISO_c, RXSM_LO_c, RXSM_SODS_c, 
        RXSM_SOE_c, stamp0_ready_dms1_c, stamp0_ready_dms2_c, 
        stamp0_ready_temp_c, stamp0_spi_miso_c, GPIO_6_M2F_c, 
        LED_HEARTBEAT_c, LED_RECORDING_c, SCLK_c, adc_clk_c, 
        adc_start_c, nCS1_c, nCS2_c, stamp0_spi_clock_c, 
        stamp0_spi_dms1_cs_c, stamp0_spi_dms2_cs_c, 
        stamp0_spi_temp_cs_c, \Memory_0.un1_APBState_1_5\, 
        mosi_cl_0, mosi_cl : std_logic;

    for all : Memory
	Use entity work.Memory(DEF_ARCH);
    for all : sb_sb
	Use entity work.sb_sb(DEF_ARCH);
    for all : STAMP
	Use entity work.STAMP(DEF_ARCH);
begin 


    stamp0_ready_dms2_ibuf : INBUF
      generic map(IOSTD => "")

      port map(PAD => stamp0_ready_dms2, Y => stamp0_ready_dms2_c);
    
    stamp0_ready_dms1_ibuf : INBUF
      generic map(IOSTD => "")

      port map(PAD => stamp0_ready_dms1, Y => stamp0_ready_dms1_c);
    
    stamp0_spi_clock_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => stamp0_spi_clock_c, PAD => stamp0_spi_clock);
    
    nCS1_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => nCS1_c, PAD => nCS1);
    
    RXSM_SODS_ibuf : INBUF
      generic map(IOSTD => "")

      port map(PAD => RXSM_SODS, Y => RXSM_SODS_c);
    
    resetn_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => NN_1, PAD => resetn);
    
    AND2_0 : AND2
      port map(A => NN_1, B => \VCC\, Y => debug_led_net_0);
    
    adc_start_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => adc_start_c, PAD => adc_start);
    
    stamp0_spi_miso_ibuf : INBUF
      generic map(IOSTD => "")

      port map(PAD => stamp0_spi_miso, Y => stamp0_spi_miso_c);
    
    MISO_ibuf : INBUF
      generic map(IOSTD => "")

      port map(PAD => MISO, Y => MISO_c);
    
    debug_led_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => \GND\, PAD => debug_led);
    
    AND2_2 : AND2
      port map(A => sb_sb_0_GPIO_3_M2F, B => \VCC\, Y => 
        adc_start_c);
    
    MOSI_obuft : TRIBUFF
      generic map(IOSTD => "")

      port map(D => mosi_1, E => mosi_cl, PAD => MOSI);
    
    AND2_0_RNIKOS1 : CLKINT
      port map(A => debug_led_net_0, Y => debug_led_net_0_arst);
    
    stamp0_spi_mosi_obuft : TRIBUFF
      generic map(IOSTD => "")

      port map(D => mosi_1_0, E => mosi_cl_0, PAD => 
        stamp0_spi_mosi);
    
    RXSM_SOE_ibuf : INBUF
      generic map(IOSTD => "")

      port map(PAD => RXSM_SOE, Y => RXSM_SOE_c);
    
    Memory_0 : Memory
      port map(sb_sb_0_STAMP_PADDR(11) => sb_sb_0_STAMP_PADDR(11), 
        sb_sb_0_STAMP_PADDR(10) => sb_sb_0_STAMP_PADDR(10), 
        sb_sb_0_STAMP_PADDR(9) => sb_sb_0_STAMP_PADDR(9), 
        sb_sb_0_STAMP_PADDR(8) => sb_sb_0_STAMP_PADDR(8), 
        sb_sb_0_STAMP_PADDR(7) => sb_sb_0_STAMP_PADDR(7), 
        sb_sb_0_STAMP_PADDR(6) => sb_sb_0_STAMP_PADDR(6), 
        sb_sb_0_STAMP_PADDR(5) => sb_sb_0_STAMP_PADDR(5), 
        sb_sb_0_STAMP_PADDR(4) => sb_sb_0_STAMP_PADDR(4), 
        sb_sb_0_STAMP_PADDR(3) => sb_sb_0_STAMP_PADDR(3), 
        sb_sb_0_STAMP_PADDR(2) => sb_sb_0_STAMP_PADDR(2), 
        sb_sb_0_STAMP_PADDR(1) => sb_sb_0_STAMP_PADDR(1), 
        sb_sb_0_STAMP_PADDR(0) => sb_sb_0_STAMP_PADDR(0), 
        dataReady_0 => \Memory_0.dataReady\(0), 
        STAMP_0_data_frame(63) => STAMP_0_data_frame(63), 
        STAMP_0_data_frame(62) => STAMP_0_data_frame(62), 
        STAMP_0_data_frame(61) => STAMP_0_data_frame(61), 
        STAMP_0_data_frame(60) => STAMP_0_data_frame(60), 
        STAMP_0_data_frame(59) => STAMP_0_data_frame(59), 
        STAMP_0_data_frame(58) => STAMP_0_data_frame(58), 
        STAMP_0_data_frame(57) => STAMP_0_data_frame(57), 
        STAMP_0_data_frame(56) => STAMP_0_data_frame(56), 
        STAMP_0_data_frame(55) => STAMP_0_data_frame(55), 
        STAMP_0_data_frame(54) => STAMP_0_data_frame(54), 
        STAMP_0_data_frame(53) => STAMP_0_data_frame(53), 
        STAMP_0_data_frame(52) => STAMP_0_data_frame(52), 
        STAMP_0_data_frame(51) => STAMP_0_data_frame(51), 
        STAMP_0_data_frame(50) => STAMP_0_data_frame(50), 
        STAMP_0_data_frame(49) => STAMP_0_data_frame(49), 
        STAMP_0_data_frame(48) => STAMP_0_data_frame(48), 
        STAMP_0_data_frame(47) => STAMP_0_data_frame(47), 
        STAMP_0_data_frame(46) => STAMP_0_data_frame(46), 
        STAMP_0_data_frame(45) => STAMP_0_data_frame(45), 
        STAMP_0_data_frame(44) => STAMP_0_data_frame(44), 
        STAMP_0_data_frame(43) => STAMP_0_data_frame(43), 
        STAMP_0_data_frame(42) => STAMP_0_data_frame(42), 
        STAMP_0_data_frame(41) => STAMP_0_data_frame(41), 
        STAMP_0_data_frame(40) => STAMP_0_data_frame(40), 
        STAMP_0_data_frame(39) => STAMP_0_data_frame(39), 
        STAMP_0_data_frame(38) => STAMP_0_data_frame(38), 
        STAMP_0_data_frame(37) => STAMP_0_data_frame(37), 
        STAMP_0_data_frame(36) => STAMP_0_data_frame(36), 
        STAMP_0_data_frame(35) => STAMP_0_data_frame(35), 
        STAMP_0_data_frame(34) => STAMP_0_data_frame(34), 
        STAMP_0_data_frame(33) => STAMP_0_data_frame(33), 
        STAMP_0_data_frame(32) => STAMP_0_data_frame(32), 
        STAMP_0_data_frame(31) => STAMP_0_data_frame(31), 
        STAMP_0_data_frame(30) => STAMP_0_data_frame(30), 
        STAMP_0_data_frame(29) => STAMP_0_data_frame(29), 
        STAMP_0_data_frame(28) => STAMP_0_data_frame(28), 
        STAMP_0_data_frame(27) => STAMP_0_data_frame(27), 
        STAMP_0_data_frame(26) => STAMP_0_data_frame(26), 
        STAMP_0_data_frame(25) => STAMP_0_data_frame(25), 
        STAMP_0_data_frame(24) => STAMP_0_data_frame(24), 
        STAMP_0_data_frame(23) => STAMP_0_data_frame(23), 
        STAMP_0_data_frame(22) => STAMP_0_data_frame(22), 
        STAMP_0_data_frame(21) => STAMP_0_data_frame(21), 
        STAMP_0_data_frame(20) => STAMP_0_data_frame(20), 
        STAMP_0_data_frame(19) => STAMP_0_data_frame(19), 
        STAMP_0_data_frame(18) => STAMP_0_data_frame(18), 
        STAMP_0_data_frame(17) => STAMP_0_data_frame(17), 
        STAMP_0_data_frame(16) => STAMP_0_data_frame(16), 
        STAMP_0_data_frame(15) => STAMP_0_data_frame(15), 
        STAMP_0_data_frame(14) => STAMP_0_data_frame(14), 
        STAMP_0_data_frame(13) => STAMP_0_data_frame(13), 
        STAMP_0_data_frame(12) => STAMP_0_data_frame(12), 
        STAMP_0_data_frame(11) => STAMP_0_data_frame(11), 
        STAMP_0_data_frame(10) => STAMP_0_data_frame(10), 
        STAMP_0_data_frame(9) => STAMP_0_data_frame(9), 
        STAMP_0_data_frame(8) => STAMP_0_data_frame(8), 
        STAMP_0_data_frame(7) => STAMP_0_data_frame(7), 
        STAMP_0_data_frame(6) => STAMP_0_data_frame(6), 
        STAMP_0_data_frame(5) => STAMP_0_data_frame(5), 
        STAMP_0_data_frame(4) => STAMP_0_data_frame(4), 
        STAMP_0_data_frame(3) => STAMP_0_data_frame(3), 
        STAMP_0_data_frame(2) => STAMP_0_data_frame(2), 
        STAMP_0_data_frame(1) => STAMP_0_data_frame(1), 
        STAMP_0_data_frame(0) => STAMP_0_data_frame(0), 
        sb_sb_0_Memory_PRDATA(31) => sb_sb_0_Memory_PRDATA(31), 
        sb_sb_0_Memory_PRDATA(30) => sb_sb_0_Memory_PRDATA(30), 
        sb_sb_0_Memory_PRDATA(29) => sb_sb_0_Memory_PRDATA(29), 
        sb_sb_0_Memory_PRDATA(28) => sb_sb_0_Memory_PRDATA(28), 
        sb_sb_0_Memory_PRDATA(27) => sb_sb_0_Memory_PRDATA(27), 
        sb_sb_0_Memory_PRDATA(26) => sb_sb_0_Memory_PRDATA(26), 
        sb_sb_0_Memory_PRDATA(25) => sb_sb_0_Memory_PRDATA(25), 
        sb_sb_0_Memory_PRDATA(24) => sb_sb_0_Memory_PRDATA(24), 
        sb_sb_0_Memory_PRDATA(23) => sb_sb_0_Memory_PRDATA(23), 
        sb_sb_0_Memory_PRDATA(22) => sb_sb_0_Memory_PRDATA(22), 
        sb_sb_0_Memory_PRDATA(21) => sb_sb_0_Memory_PRDATA(21), 
        sb_sb_0_Memory_PRDATA(20) => sb_sb_0_Memory_PRDATA(20), 
        sb_sb_0_Memory_PRDATA(19) => sb_sb_0_Memory_PRDATA(19), 
        sb_sb_0_Memory_PRDATA(18) => sb_sb_0_Memory_PRDATA(18), 
        sb_sb_0_Memory_PRDATA(17) => sb_sb_0_Memory_PRDATA(17), 
        sb_sb_0_Memory_PRDATA(16) => sb_sb_0_Memory_PRDATA(16), 
        sb_sb_0_Memory_PRDATA(15) => sb_sb_0_Memory_PRDATA(15), 
        sb_sb_0_Memory_PRDATA(14) => sb_sb_0_Memory_PRDATA(14), 
        sb_sb_0_Memory_PRDATA(13) => sb_sb_0_Memory_PRDATA(13), 
        sb_sb_0_Memory_PRDATA(12) => sb_sb_0_Memory_PRDATA(12), 
        sb_sb_0_Memory_PRDATA(11) => sb_sb_0_Memory_PRDATA(11), 
        sb_sb_0_Memory_PRDATA(10) => sb_sb_0_Memory_PRDATA(10), 
        sb_sb_0_Memory_PRDATA(9) => sb_sb_0_Memory_PRDATA(9), 
        sb_sb_0_Memory_PRDATA(8) => sb_sb_0_Memory_PRDATA(8), 
        sb_sb_0_Memory_PRDATA(7) => sb_sb_0_Memory_PRDATA(7), 
        sb_sb_0_Memory_PRDATA(6) => sb_sb_0_Memory_PRDATA(6), 
        sb_sb_0_Memory_PRDATA(5) => sb_sb_0_Memory_PRDATA(5), 
        sb_sb_0_Memory_PRDATA(4) => sb_sb_0_Memory_PRDATA(4), 
        sb_sb_0_Memory_PRDATA(3) => sb_sb_0_Memory_PRDATA(3), 
        sb_sb_0_Memory_PRDATA(2) => sb_sb_0_Memory_PRDATA(2), 
        sb_sb_0_Memory_PRDATA(1) => sb_sb_0_Memory_PRDATA(1), 
        sb_sb_0_Memory_PRDATA(0) => sb_sb_0_Memory_PRDATA(0), 
        sb_sb_0_STAMP_PWDATA(31) => sb_sb_0_STAMP_PWDATA(31), 
        sb_sb_0_STAMP_PWDATA(30) => sb_sb_0_STAMP_PWDATA(30), 
        sb_sb_0_STAMP_PWDATA(29) => sb_sb_0_STAMP_PWDATA(29), 
        sb_sb_0_STAMP_PWDATA(28) => sb_sb_0_STAMP_PWDATA(28), 
        sb_sb_0_STAMP_PWDATA(27) => sb_sb_0_STAMP_PWDATA(27), 
        sb_sb_0_STAMP_PWDATA(26) => sb_sb_0_STAMP_PWDATA(26), 
        sb_sb_0_STAMP_PWDATA(25) => sb_sb_0_STAMP_PWDATA(25), 
        sb_sb_0_STAMP_PWDATA(24) => sb_sb_0_STAMP_PWDATA(24), 
        sb_sb_0_STAMP_PWDATA(23) => sb_sb_0_STAMP_PWDATA(23), 
        sb_sb_0_STAMP_PWDATA(22) => sb_sb_0_STAMP_PWDATA(22), 
        sb_sb_0_STAMP_PWDATA(21) => sb_sb_0_STAMP_PWDATA(21), 
        sb_sb_0_STAMP_PWDATA(20) => sb_sb_0_STAMP_PWDATA(20), 
        sb_sb_0_STAMP_PWDATA(19) => sb_sb_0_STAMP_PWDATA(19), 
        sb_sb_0_STAMP_PWDATA(18) => sb_sb_0_STAMP_PWDATA(18), 
        sb_sb_0_STAMP_PWDATA(17) => sb_sb_0_STAMP_PWDATA(17), 
        sb_sb_0_STAMP_PWDATA(16) => sb_sb_0_STAMP_PWDATA(16), 
        sb_sb_0_STAMP_PWDATA(15) => sb_sb_0_STAMP_PWDATA(15), 
        sb_sb_0_STAMP_PWDATA(14) => sb_sb_0_STAMP_PWDATA(14), 
        sb_sb_0_STAMP_PWDATA(13) => sb_sb_0_STAMP_PWDATA(13), 
        sb_sb_0_STAMP_PWDATA(12) => sb_sb_0_STAMP_PWDATA(12), 
        sb_sb_0_STAMP_PWDATA(11) => sb_sb_0_STAMP_PWDATA(11), 
        sb_sb_0_STAMP_PWDATA(10) => sb_sb_0_STAMP_PWDATA(10), 
        sb_sb_0_STAMP_PWDATA(9) => sb_sb_0_STAMP_PWDATA(9), 
        sb_sb_0_STAMP_PWDATA(8) => sb_sb_0_STAMP_PWDATA(8), 
        sb_sb_0_STAMP_PWDATA(7) => sb_sb_0_STAMP_PWDATA(7), 
        sb_sb_0_STAMP_PWDATA(6) => sb_sb_0_STAMP_PWDATA(6), 
        sb_sb_0_STAMP_PWDATA(5) => sb_sb_0_STAMP_PWDATA(5), 
        sb_sb_0_STAMP_PWDATA(4) => sb_sb_0_STAMP_PWDATA(4), 
        sb_sb_0_STAMP_PWDATA(3) => sb_sb_0_STAMP_PWDATA(3), 
        sb_sb_0_STAMP_PWDATA(2) => sb_sb_0_STAMP_PWDATA(2), 
        sb_sb_0_STAMP_PWDATA(1) => sb_sb_0_STAMP_PWDATA(1), 
        sb_sb_0_STAMP_PWDATA(0) => sb_sb_0_STAMP_PWDATA(0), 
        nCS1_c => nCS1_c, nCS2_c => nCS2_c, MISO_c => MISO_c, 
        SCLK_c => SCLK_c, mosi_1 => mosi_1, mosi_cl => mosi_cl, 
        sb_sb_0_STAMP_PENABLE => sb_sb_0_STAMP_PENABLE, 
        sb_sb_0_STAMP_PWRITE => sb_sb_0_STAMP_PWRITE, 
        sb_sb_0_Memory_PSELx => sb_sb_0_Memory_PSELx, 
        un1_APBState_1_5_1z => \Memory_0.un1_APBState_1_5\, 
        resetn => NN_1, sb_sb_0_Memory_PREADY => 
        sb_sb_0_Memory_PREADY, GPIO_6_M2F_c => GPIO_6_M2F_c, 
        sb_sb_0_FIC_0_CLK => sb_sb_0_FIC_0_CLK, resetn_arst => 
        resetn_arst);
    
    sb_sb_0 : sb_sb
      port map(sb_sb_0_STAMP_PADDR(11) => sb_sb_0_STAMP_PADDR(11), 
        sb_sb_0_STAMP_PADDR(10) => sb_sb_0_STAMP_PADDR(10), 
        sb_sb_0_STAMP_PADDR(9) => sb_sb_0_STAMP_PADDR(9), 
        sb_sb_0_STAMP_PADDR(8) => sb_sb_0_STAMP_PADDR(8), 
        sb_sb_0_STAMP_PADDR(7) => sb_sb_0_STAMP_PADDR(7), 
        sb_sb_0_STAMP_PADDR(6) => sb_sb_0_STAMP_PADDR(6), 
        sb_sb_0_STAMP_PADDR(5) => sb_sb_0_STAMP_PADDR(5), 
        sb_sb_0_STAMP_PADDR(4) => sb_sb_0_STAMP_PADDR(4), 
        sb_sb_0_STAMP_PADDR(3) => sb_sb_0_STAMP_PADDR(3), 
        sb_sb_0_STAMP_PADDR(2) => sb_sb_0_STAMP_PADDR(2), 
        sb_sb_0_STAMP_PADDR(1) => sb_sb_0_STAMP_PADDR(1), 
        sb_sb_0_STAMP_PADDR(0) => sb_sb_0_STAMP_PADDR(0), 
        sb_sb_0_STAMP_PWDATA(31) => sb_sb_0_STAMP_PWDATA(31), 
        sb_sb_0_STAMP_PWDATA(30) => sb_sb_0_STAMP_PWDATA(30), 
        sb_sb_0_STAMP_PWDATA(29) => sb_sb_0_STAMP_PWDATA(29), 
        sb_sb_0_STAMP_PWDATA(28) => sb_sb_0_STAMP_PWDATA(28), 
        sb_sb_0_STAMP_PWDATA(27) => sb_sb_0_STAMP_PWDATA(27), 
        sb_sb_0_STAMP_PWDATA(26) => sb_sb_0_STAMP_PWDATA(26), 
        sb_sb_0_STAMP_PWDATA(25) => sb_sb_0_STAMP_PWDATA(25), 
        sb_sb_0_STAMP_PWDATA(24) => sb_sb_0_STAMP_PWDATA(24), 
        sb_sb_0_STAMP_PWDATA(23) => sb_sb_0_STAMP_PWDATA(23), 
        sb_sb_0_STAMP_PWDATA(22) => sb_sb_0_STAMP_PWDATA(22), 
        sb_sb_0_STAMP_PWDATA(21) => sb_sb_0_STAMP_PWDATA(21), 
        sb_sb_0_STAMP_PWDATA(20) => sb_sb_0_STAMP_PWDATA(20), 
        sb_sb_0_STAMP_PWDATA(19) => sb_sb_0_STAMP_PWDATA(19), 
        sb_sb_0_STAMP_PWDATA(18) => sb_sb_0_STAMP_PWDATA(18), 
        sb_sb_0_STAMP_PWDATA(17) => sb_sb_0_STAMP_PWDATA(17), 
        sb_sb_0_STAMP_PWDATA(16) => sb_sb_0_STAMP_PWDATA(16), 
        sb_sb_0_STAMP_PWDATA(15) => sb_sb_0_STAMP_PWDATA(15), 
        sb_sb_0_STAMP_PWDATA(14) => sb_sb_0_STAMP_PWDATA(14), 
        sb_sb_0_STAMP_PWDATA(13) => sb_sb_0_STAMP_PWDATA(13), 
        sb_sb_0_STAMP_PWDATA(12) => sb_sb_0_STAMP_PWDATA(12), 
        sb_sb_0_STAMP_PWDATA(11) => sb_sb_0_STAMP_PWDATA(11), 
        sb_sb_0_STAMP_PWDATA(10) => sb_sb_0_STAMP_PWDATA(10), 
        sb_sb_0_STAMP_PWDATA(9) => sb_sb_0_STAMP_PWDATA(9), 
        sb_sb_0_STAMP_PWDATA(8) => sb_sb_0_STAMP_PWDATA(8), 
        sb_sb_0_STAMP_PWDATA(7) => sb_sb_0_STAMP_PWDATA(7), 
        sb_sb_0_STAMP_PWDATA(6) => sb_sb_0_STAMP_PWDATA(6), 
        sb_sb_0_STAMP_PWDATA(5) => sb_sb_0_STAMP_PWDATA(5), 
        sb_sb_0_STAMP_PWDATA(4) => sb_sb_0_STAMP_PWDATA(4), 
        sb_sb_0_STAMP_PWDATA(3) => sb_sb_0_STAMP_PWDATA(3), 
        sb_sb_0_STAMP_PWDATA(2) => sb_sb_0_STAMP_PWDATA(2), 
        sb_sb_0_STAMP_PWDATA(1) => sb_sb_0_STAMP_PWDATA(1), 
        sb_sb_0_STAMP_PWDATA(0) => sb_sb_0_STAMP_PWDATA(0), 
        dataReady_0 => \Memory_0.dataReady\(0), 
        sb_sb_0_Memory_PRDATA(31) => sb_sb_0_Memory_PRDATA(31), 
        sb_sb_0_Memory_PRDATA(30) => sb_sb_0_Memory_PRDATA(30), 
        sb_sb_0_Memory_PRDATA(29) => sb_sb_0_Memory_PRDATA(29), 
        sb_sb_0_Memory_PRDATA(28) => sb_sb_0_Memory_PRDATA(28), 
        sb_sb_0_Memory_PRDATA(27) => sb_sb_0_Memory_PRDATA(27), 
        sb_sb_0_Memory_PRDATA(26) => sb_sb_0_Memory_PRDATA(26), 
        sb_sb_0_Memory_PRDATA(25) => sb_sb_0_Memory_PRDATA(25), 
        sb_sb_0_Memory_PRDATA(24) => sb_sb_0_Memory_PRDATA(24), 
        sb_sb_0_Memory_PRDATA(23) => sb_sb_0_Memory_PRDATA(23), 
        sb_sb_0_Memory_PRDATA(22) => sb_sb_0_Memory_PRDATA(22), 
        sb_sb_0_Memory_PRDATA(21) => sb_sb_0_Memory_PRDATA(21), 
        sb_sb_0_Memory_PRDATA(20) => sb_sb_0_Memory_PRDATA(20), 
        sb_sb_0_Memory_PRDATA(19) => sb_sb_0_Memory_PRDATA(19), 
        sb_sb_0_Memory_PRDATA(18) => sb_sb_0_Memory_PRDATA(18), 
        sb_sb_0_Memory_PRDATA(17) => sb_sb_0_Memory_PRDATA(17), 
        sb_sb_0_Memory_PRDATA(16) => sb_sb_0_Memory_PRDATA(16), 
        sb_sb_0_Memory_PRDATA(15) => sb_sb_0_Memory_PRDATA(15), 
        sb_sb_0_Memory_PRDATA(14) => sb_sb_0_Memory_PRDATA(14), 
        sb_sb_0_Memory_PRDATA(13) => sb_sb_0_Memory_PRDATA(13), 
        sb_sb_0_Memory_PRDATA(12) => sb_sb_0_Memory_PRDATA(12), 
        sb_sb_0_Memory_PRDATA(11) => sb_sb_0_Memory_PRDATA(11), 
        sb_sb_0_Memory_PRDATA(10) => sb_sb_0_Memory_PRDATA(10), 
        sb_sb_0_Memory_PRDATA(9) => sb_sb_0_Memory_PRDATA(9), 
        sb_sb_0_Memory_PRDATA(8) => sb_sb_0_Memory_PRDATA(8), 
        sb_sb_0_Memory_PRDATA(7) => sb_sb_0_Memory_PRDATA(7), 
        sb_sb_0_Memory_PRDATA(6) => sb_sb_0_Memory_PRDATA(6), 
        sb_sb_0_Memory_PRDATA(5) => sb_sb_0_Memory_PRDATA(5), 
        sb_sb_0_Memory_PRDATA(4) => sb_sb_0_Memory_PRDATA(4), 
        sb_sb_0_Memory_PRDATA(3) => sb_sb_0_Memory_PRDATA(3), 
        sb_sb_0_Memory_PRDATA(2) => sb_sb_0_Memory_PRDATA(2), 
        sb_sb_0_Memory_PRDATA(1) => sb_sb_0_Memory_PRDATA(1), 
        sb_sb_0_Memory_PRDATA(0) => sb_sb_0_Memory_PRDATA(0), 
        sb_sb_0_STAMP_PRDATA(31) => sb_sb_0_STAMP_PRDATA(31), 
        sb_sb_0_STAMP_PRDATA(30) => sb_sb_0_STAMP_PRDATA(30), 
        sb_sb_0_STAMP_PRDATA(29) => sb_sb_0_STAMP_PRDATA(29), 
        sb_sb_0_STAMP_PRDATA(28) => sb_sb_0_STAMP_PRDATA(28), 
        sb_sb_0_STAMP_PRDATA(27) => sb_sb_0_STAMP_PRDATA(27), 
        sb_sb_0_STAMP_PRDATA(26) => sb_sb_0_STAMP_PRDATA(26), 
        sb_sb_0_STAMP_PRDATA(25) => sb_sb_0_STAMP_PRDATA(25), 
        sb_sb_0_STAMP_PRDATA(24) => sb_sb_0_STAMP_PRDATA(24), 
        sb_sb_0_STAMP_PRDATA(23) => sb_sb_0_STAMP_PRDATA(23), 
        sb_sb_0_STAMP_PRDATA(22) => sb_sb_0_STAMP_PRDATA(22), 
        sb_sb_0_STAMP_PRDATA(21) => sb_sb_0_STAMP_PRDATA(21), 
        sb_sb_0_STAMP_PRDATA(20) => sb_sb_0_STAMP_PRDATA(20), 
        sb_sb_0_STAMP_PRDATA(19) => sb_sb_0_STAMP_PRDATA(19), 
        sb_sb_0_STAMP_PRDATA(18) => sb_sb_0_STAMP_PRDATA(18), 
        sb_sb_0_STAMP_PRDATA(17) => sb_sb_0_STAMP_PRDATA(17), 
        sb_sb_0_STAMP_PRDATA(16) => sb_sb_0_STAMP_PRDATA(16), 
        sb_sb_0_STAMP_PRDATA(15) => sb_sb_0_STAMP_PRDATA(15), 
        sb_sb_0_STAMP_PRDATA(14) => sb_sb_0_STAMP_PRDATA(14), 
        sb_sb_0_STAMP_PRDATA(13) => sb_sb_0_STAMP_PRDATA(13), 
        sb_sb_0_STAMP_PRDATA(12) => sb_sb_0_STAMP_PRDATA(12), 
        sb_sb_0_STAMP_PRDATA(11) => sb_sb_0_STAMP_PRDATA(11), 
        sb_sb_0_STAMP_PRDATA(10) => sb_sb_0_STAMP_PRDATA(10), 
        sb_sb_0_STAMP_PRDATA(9) => sb_sb_0_STAMP_PRDATA(9), 
        sb_sb_0_STAMP_PRDATA(8) => sb_sb_0_STAMP_PRDATA(8), 
        sb_sb_0_STAMP_PRDATA(7) => sb_sb_0_STAMP_PRDATA(7), 
        sb_sb_0_STAMP_PRDATA(6) => sb_sb_0_STAMP_PRDATA(6), 
        sb_sb_0_STAMP_PRDATA(5) => sb_sb_0_STAMP_PRDATA(5), 
        sb_sb_0_STAMP_PRDATA(4) => sb_sb_0_STAMP_PRDATA(4), 
        sb_sb_0_STAMP_PRDATA(3) => sb_sb_0_STAMP_PRDATA(3), 
        sb_sb_0_STAMP_PRDATA(2) => sb_sb_0_STAMP_PRDATA(2), 
        sb_sb_0_STAMP_PRDATA(1) => sb_sb_0_STAMP_PRDATA(1), 
        sb_sb_0_STAMP_PRDATA(0) => sb_sb_0_STAMP_PRDATA(0), TM_TX
         => TM_TX, TM_RX => TM_RX, DAPI_TX => DAPI_TX, DAPI_RX
         => DAPI_RX, sb_sb_0_GPIO_3_M2F => sb_sb_0_GPIO_3_M2F, 
        sb_sb_0_GPIO_4_M2F => sb_sb_0_GPIO_4_M2F, 
        sb_sb_0_STAMP_PENABLE => sb_sb_0_STAMP_PENABLE, 
        sb_sb_0_STAMP_PWRITE => sb_sb_0_STAMP_PWRITE, 
        LED_HEARTBEAT_c => LED_HEARTBEAT_c, LED_RECORDING_c => 
        LED_RECORDING_c, GPIO_6_M2F_c => GPIO_6_M2F_c, RXSM_LO_c
         => RXSM_LO_c, RXSM_SOE_c => RXSM_SOE_c, RXSM_SODS_c => 
        RXSM_SODS_c, sb_sb_0_Memory_PSELx => sb_sb_0_Memory_PSELx, 
        sb_sb_0_STAMP_PSELx => sb_sb_0_STAMP_PSELx, 
        sb_sb_0_Memory_PREADY => sb_sb_0_Memory_PREADY, 
        sb_sb_0_STAMP_PREADY => sb_sb_0_STAMP_PREADY, 
        sb_sb_0_FIC_0_CLK => sb_sb_0_FIC_0_CLK, adc_clk_c => 
        adc_clk_c, DEVRST_N => DEVRST_N, sb_sb_0_POWER_ON_RESET_N
         => sb_sb_0_POWER_ON_RESET_N);
    
    ResetAND_RNIMHJB : CLKINT
      port map(A => NN_1, Y => resetn_arst);
    
    stamp0_spi_dms2_cs_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => stamp0_spi_dms2_cs_c, PAD => 
        stamp0_spi_dms2_cs);
    
    STAMP_0 : STAMP
      port map(sb_sb_0_STAMP_PADDR(11) => sb_sb_0_STAMP_PADDR(11), 
        sb_sb_0_STAMP_PADDR(10) => sb_sb_0_STAMP_PADDR(10), 
        sb_sb_0_STAMP_PADDR(9) => sb_sb_0_STAMP_PADDR(9), 
        sb_sb_0_STAMP_PADDR(8) => sb_sb_0_STAMP_PADDR(8), 
        sb_sb_0_STAMP_PADDR(7) => sb_sb_0_STAMP_PADDR(7), 
        sb_sb_0_STAMP_PADDR(6) => sb_sb_0_STAMP_PADDR(6), 
        sb_sb_0_STAMP_PADDR(5) => sb_sb_0_STAMP_PADDR(5), 
        sb_sb_0_STAMP_PADDR(4) => sb_sb_0_STAMP_PADDR(4), 
        sb_sb_0_STAMP_PADDR(3) => sb_sb_0_STAMP_PADDR(3), 
        sb_sb_0_STAMP_PADDR(2) => sb_sb_0_STAMP_PADDR(2), 
        STAMP_0_data_frame(63) => STAMP_0_data_frame(63), 
        STAMP_0_data_frame(62) => STAMP_0_data_frame(62), 
        STAMP_0_data_frame(61) => STAMP_0_data_frame(61), 
        STAMP_0_data_frame(60) => STAMP_0_data_frame(60), 
        STAMP_0_data_frame(59) => STAMP_0_data_frame(59), 
        STAMP_0_data_frame(58) => STAMP_0_data_frame(58), 
        STAMP_0_data_frame(57) => STAMP_0_data_frame(57), 
        STAMP_0_data_frame(56) => STAMP_0_data_frame(56), 
        STAMP_0_data_frame(55) => STAMP_0_data_frame(55), 
        STAMP_0_data_frame(54) => STAMP_0_data_frame(54), 
        STAMP_0_data_frame(53) => STAMP_0_data_frame(53), 
        STAMP_0_data_frame(52) => STAMP_0_data_frame(52), 
        STAMP_0_data_frame(51) => STAMP_0_data_frame(51), 
        STAMP_0_data_frame(50) => STAMP_0_data_frame(50), 
        STAMP_0_data_frame(49) => STAMP_0_data_frame(49), 
        STAMP_0_data_frame(48) => STAMP_0_data_frame(48), 
        STAMP_0_data_frame(47) => STAMP_0_data_frame(47), 
        STAMP_0_data_frame(46) => STAMP_0_data_frame(46), 
        STAMP_0_data_frame(45) => STAMP_0_data_frame(45), 
        STAMP_0_data_frame(44) => STAMP_0_data_frame(44), 
        STAMP_0_data_frame(43) => STAMP_0_data_frame(43), 
        STAMP_0_data_frame(42) => STAMP_0_data_frame(42), 
        STAMP_0_data_frame(41) => STAMP_0_data_frame(41), 
        STAMP_0_data_frame(40) => STAMP_0_data_frame(40), 
        STAMP_0_data_frame(39) => STAMP_0_data_frame(39), 
        STAMP_0_data_frame(38) => STAMP_0_data_frame(38), 
        STAMP_0_data_frame(37) => STAMP_0_data_frame(37), 
        STAMP_0_data_frame(36) => STAMP_0_data_frame(36), 
        STAMP_0_data_frame(35) => STAMP_0_data_frame(35), 
        STAMP_0_data_frame(34) => STAMP_0_data_frame(34), 
        STAMP_0_data_frame(33) => STAMP_0_data_frame(33), 
        STAMP_0_data_frame(32) => STAMP_0_data_frame(32), 
        STAMP_0_data_frame(31) => STAMP_0_data_frame(31), 
        STAMP_0_data_frame(30) => STAMP_0_data_frame(30), 
        STAMP_0_data_frame(29) => STAMP_0_data_frame(29), 
        STAMP_0_data_frame(28) => STAMP_0_data_frame(28), 
        STAMP_0_data_frame(27) => STAMP_0_data_frame(27), 
        STAMP_0_data_frame(26) => STAMP_0_data_frame(26), 
        STAMP_0_data_frame(25) => STAMP_0_data_frame(25), 
        STAMP_0_data_frame(24) => STAMP_0_data_frame(24), 
        STAMP_0_data_frame(23) => STAMP_0_data_frame(23), 
        STAMP_0_data_frame(22) => STAMP_0_data_frame(22), 
        STAMP_0_data_frame(21) => STAMP_0_data_frame(21), 
        STAMP_0_data_frame(20) => STAMP_0_data_frame(20), 
        STAMP_0_data_frame(19) => STAMP_0_data_frame(19), 
        STAMP_0_data_frame(18) => STAMP_0_data_frame(18), 
        STAMP_0_data_frame(17) => STAMP_0_data_frame(17), 
        STAMP_0_data_frame(16) => STAMP_0_data_frame(16), 
        STAMP_0_data_frame(15) => STAMP_0_data_frame(15), 
        STAMP_0_data_frame(14) => STAMP_0_data_frame(14), 
        STAMP_0_data_frame(13) => STAMP_0_data_frame(13), 
        STAMP_0_data_frame(12) => STAMP_0_data_frame(12), 
        STAMP_0_data_frame(11) => STAMP_0_data_frame(11), 
        STAMP_0_data_frame(10) => STAMP_0_data_frame(10), 
        STAMP_0_data_frame(9) => STAMP_0_data_frame(9), 
        STAMP_0_data_frame(8) => STAMP_0_data_frame(8), 
        STAMP_0_data_frame(7) => STAMP_0_data_frame(7), 
        STAMP_0_data_frame(6) => STAMP_0_data_frame(6), 
        STAMP_0_data_frame(5) => STAMP_0_data_frame(5), 
        STAMP_0_data_frame(4) => STAMP_0_data_frame(4), 
        STAMP_0_data_frame(3) => STAMP_0_data_frame(3), 
        STAMP_0_data_frame(2) => STAMP_0_data_frame(2), 
        STAMP_0_data_frame(1) => STAMP_0_data_frame(1), 
        STAMP_0_data_frame(0) => STAMP_0_data_frame(0), 
        sb_sb_0_STAMP_PRDATA(31) => sb_sb_0_STAMP_PRDATA(31), 
        sb_sb_0_STAMP_PRDATA(30) => sb_sb_0_STAMP_PRDATA(30), 
        sb_sb_0_STAMP_PRDATA(29) => sb_sb_0_STAMP_PRDATA(29), 
        sb_sb_0_STAMP_PRDATA(28) => sb_sb_0_STAMP_PRDATA(28), 
        sb_sb_0_STAMP_PRDATA(27) => sb_sb_0_STAMP_PRDATA(27), 
        sb_sb_0_STAMP_PRDATA(26) => sb_sb_0_STAMP_PRDATA(26), 
        sb_sb_0_STAMP_PRDATA(25) => sb_sb_0_STAMP_PRDATA(25), 
        sb_sb_0_STAMP_PRDATA(24) => sb_sb_0_STAMP_PRDATA(24), 
        sb_sb_0_STAMP_PRDATA(23) => sb_sb_0_STAMP_PRDATA(23), 
        sb_sb_0_STAMP_PRDATA(22) => sb_sb_0_STAMP_PRDATA(22), 
        sb_sb_0_STAMP_PRDATA(21) => sb_sb_0_STAMP_PRDATA(21), 
        sb_sb_0_STAMP_PRDATA(20) => sb_sb_0_STAMP_PRDATA(20), 
        sb_sb_0_STAMP_PRDATA(19) => sb_sb_0_STAMP_PRDATA(19), 
        sb_sb_0_STAMP_PRDATA(18) => sb_sb_0_STAMP_PRDATA(18), 
        sb_sb_0_STAMP_PRDATA(17) => sb_sb_0_STAMP_PRDATA(17), 
        sb_sb_0_STAMP_PRDATA(16) => sb_sb_0_STAMP_PRDATA(16), 
        sb_sb_0_STAMP_PRDATA(15) => sb_sb_0_STAMP_PRDATA(15), 
        sb_sb_0_STAMP_PRDATA(14) => sb_sb_0_STAMP_PRDATA(14), 
        sb_sb_0_STAMP_PRDATA(13) => sb_sb_0_STAMP_PRDATA(13), 
        sb_sb_0_STAMP_PRDATA(12) => sb_sb_0_STAMP_PRDATA(12), 
        sb_sb_0_STAMP_PRDATA(11) => sb_sb_0_STAMP_PRDATA(11), 
        sb_sb_0_STAMP_PRDATA(10) => sb_sb_0_STAMP_PRDATA(10), 
        sb_sb_0_STAMP_PRDATA(9) => sb_sb_0_STAMP_PRDATA(9), 
        sb_sb_0_STAMP_PRDATA(8) => sb_sb_0_STAMP_PRDATA(8), 
        sb_sb_0_STAMP_PRDATA(7) => sb_sb_0_STAMP_PRDATA(7), 
        sb_sb_0_STAMP_PRDATA(6) => sb_sb_0_STAMP_PRDATA(6), 
        sb_sb_0_STAMP_PRDATA(5) => sb_sb_0_STAMP_PRDATA(5), 
        sb_sb_0_STAMP_PRDATA(4) => sb_sb_0_STAMP_PRDATA(4), 
        sb_sb_0_STAMP_PRDATA(3) => sb_sb_0_STAMP_PRDATA(3), 
        sb_sb_0_STAMP_PRDATA(2) => sb_sb_0_STAMP_PRDATA(2), 
        sb_sb_0_STAMP_PRDATA(1) => sb_sb_0_STAMP_PRDATA(1), 
        sb_sb_0_STAMP_PRDATA(0) => sb_sb_0_STAMP_PRDATA(0), 
        dataReady_0 => \Memory_0.dataReady\(0), 
        sb_sb_0_STAMP_PWDATA(31) => sb_sb_0_STAMP_PWDATA(31), 
        sb_sb_0_STAMP_PWDATA(30) => sb_sb_0_STAMP_PWDATA(30), 
        sb_sb_0_STAMP_PWDATA(29) => sb_sb_0_STAMP_PWDATA(29), 
        sb_sb_0_STAMP_PWDATA(28) => sb_sb_0_STAMP_PWDATA(28), 
        sb_sb_0_STAMP_PWDATA(27) => sb_sb_0_STAMP_PWDATA(27), 
        sb_sb_0_STAMP_PWDATA(26) => sb_sb_0_STAMP_PWDATA(26), 
        sb_sb_0_STAMP_PWDATA(25) => sb_sb_0_STAMP_PWDATA(25), 
        sb_sb_0_STAMP_PWDATA(24) => sb_sb_0_STAMP_PWDATA(24), 
        sb_sb_0_STAMP_PWDATA(23) => sb_sb_0_STAMP_PWDATA(23), 
        sb_sb_0_STAMP_PWDATA(22) => sb_sb_0_STAMP_PWDATA(22), 
        sb_sb_0_STAMP_PWDATA(21) => sb_sb_0_STAMP_PWDATA(21), 
        sb_sb_0_STAMP_PWDATA(20) => sb_sb_0_STAMP_PWDATA(20), 
        sb_sb_0_STAMP_PWDATA(19) => sb_sb_0_STAMP_PWDATA(19), 
        sb_sb_0_STAMP_PWDATA(18) => sb_sb_0_STAMP_PWDATA(18), 
        sb_sb_0_STAMP_PWDATA(17) => sb_sb_0_STAMP_PWDATA(17), 
        sb_sb_0_STAMP_PWDATA(16) => sb_sb_0_STAMP_PWDATA(16), 
        sb_sb_0_STAMP_PWDATA(15) => sb_sb_0_STAMP_PWDATA(15), 
        sb_sb_0_STAMP_PWDATA(14) => sb_sb_0_STAMP_PWDATA(14), 
        sb_sb_0_STAMP_PWDATA(13) => sb_sb_0_STAMP_PWDATA(13), 
        sb_sb_0_STAMP_PWDATA(12) => sb_sb_0_STAMP_PWDATA(12), 
        sb_sb_0_STAMP_PWDATA(11) => sb_sb_0_STAMP_PWDATA(11), 
        sb_sb_0_STAMP_PWDATA(10) => sb_sb_0_STAMP_PWDATA(10), 
        sb_sb_0_STAMP_PWDATA(9) => sb_sb_0_STAMP_PWDATA(9), 
        sb_sb_0_STAMP_PWDATA(8) => sb_sb_0_STAMP_PWDATA(8), 
        sb_sb_0_STAMP_PWDATA(7) => sb_sb_0_STAMP_PWDATA(7), 
        sb_sb_0_STAMP_PWDATA(6) => sb_sb_0_STAMP_PWDATA(6), 
        sb_sb_0_STAMP_PWDATA(5) => sb_sb_0_STAMP_PWDATA(5), 
        sb_sb_0_STAMP_PWDATA(4) => sb_sb_0_STAMP_PWDATA(4), 
        sb_sb_0_STAMP_PWDATA(3) => sb_sb_0_STAMP_PWDATA(3), 
        sb_sb_0_STAMP_PWDATA(2) => sb_sb_0_STAMP_PWDATA(2), 
        sb_sb_0_STAMP_PWDATA(1) => sb_sb_0_STAMP_PWDATA(1), 
        sb_sb_0_STAMP_PWDATA(0) => sb_sb_0_STAMP_PWDATA(0), 
        stamp0_spi_miso_c => stamp0_spi_miso_c, 
        stamp0_spi_clock_c => stamp0_spi_clock_c, mosi_1_0 => 
        mosi_1_0, mosi_cl_0 => mosi_cl_0, sb_sb_0_STAMP_PSELx => 
        sb_sb_0_STAMP_PSELx, sb_sb_0_STAMP_PENABLE => 
        sb_sb_0_STAMP_PENABLE, un1_APBState_1_5 => 
        \Memory_0.un1_APBState_1_5\, sb_sb_0_STAMP_PWRITE => 
        sb_sb_0_STAMP_PWRITE, sb_sb_0_STAMP_PREADY => 
        sb_sb_0_STAMP_PREADY, debug_led_net_0 => debug_led_net_0, 
        stamp0_spi_dms1_cs_c => stamp0_spi_dms1_cs_c, 
        stamp0_spi_temp_cs_c => stamp0_spi_temp_cs_c, 
        stamp0_spi_dms2_cs_c => stamp0_spi_dms2_cs_c, 
        sb_sb_0_FIC_0_CLK => sb_sb_0_FIC_0_CLK, 
        debug_led_net_0_arst => debug_led_net_0_arst, 
        stamp0_ready_dms1_c => stamp0_ready_dms1_c, 
        stamp0_ready_temp_c => stamp0_ready_temp_c, 
        stamp0_ready_dms2_c => stamp0_ready_dms2_c);
    
    stamp0_ready_temp_ibuf : INBUF
      generic map(IOSTD => "")

      port map(PAD => stamp0_ready_temp, Y => stamp0_ready_temp_c);
    
    GPIO_6_M2F_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => GPIO_6_M2F_c, PAD => GPIO_6_M2F);
    
    LED_HEARTBEAT_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => LED_HEARTBEAT_c, PAD => LED_HEARTBEAT);
    
    SCLK_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => SCLK_c, PAD => SCLK);
    
    GND_Z : GND
      port map(Y => \GND\);
    
    VCC_Z : VCC
      port map(Y => \VCC\);
    
    adc_clk_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => adc_clk_c, PAD => adc_clk);
    
    stamp0_spi_temp_cs_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => stamp0_spi_temp_cs_c, PAD => 
        stamp0_spi_temp_cs);
    
    ResetAND : AND2
      port map(A => sb_sb_0_POWER_ON_RESET_N, B => 
        sb_sb_0_GPIO_4_M2F, Y => NN_1);
    
    LED_RECORDING_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => LED_RECORDING_c, PAD => LED_RECORDING);
    
    nCS2_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => nCS2_c, PAD => nCS2);
    
    RXSM_LO_ibuf : INBUF
      generic map(IOSTD => "")

      port map(PAD => RXSM_LO, Y => RXSM_LO_c);
    
    stamp0_spi_dms1_cs_obuf : OUTBUF
      generic map(IOSTD => "")

      port map(D => stamp0_spi_dms1_cs_c, PAD => 
        stamp0_spi_dms1_cs);
    

end DEF_ARCH; 
